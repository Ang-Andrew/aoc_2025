localparam N = 496;
localparam N_PADDED = 496;
localparam DEPTH = 124;
