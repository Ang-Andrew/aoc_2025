localparam MAX_ROWS = 32;
localparam STREAM_DEPTH = 1312;
