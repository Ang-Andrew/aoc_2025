localparam NUM_RANGES = 174;
localparam NUM_IDS = 1000;
