localparam WIDTH = 3724;
localparam HEIGHT = 5;
localparam MEM_SIZE = 18620;
