// Day 3 ROM: 200 precomputed line scores
// Total sum: 17092
module rom_hardcoded (
    input wire [7:0] addr,
    output reg [31:0] data
);

    always @(*) begin
        case(addr)
            8'd0: data = 32'h0000004c;
            8'd1: data = 32'h00000063;
            8'd2: data = 32'h0000005e;
            8'd3: data = 32'h00000062;
            8'd4: data = 32'h00000058;
            8'd5: data = 32'h00000063;
            8'd6: data = 32'h00000063;
            8'd7: data = 32'h00000063;
            8'd8: data = 32'h00000062;
            8'd9: data = 32'h00000062;
            8'd10: data = 32'h00000058;
            8'd11: data = 32'h00000062;
            8'd12: data = 32'h00000063;
            8'd13: data = 32'h00000042;
            8'd14: data = 32'h00000058;
            8'd15: data = 32'h00000061;
            8'd16: data = 32'h00000063;
            8'd17: data = 32'h00000058;
            8'd18: data = 32'h00000060;
            8'd19: data = 32'h00000058;
            8'd20: data = 32'h00000060;
            8'd21: data = 32'h00000062;
            8'd22: data = 32'h00000063;
            8'd23: data = 32'h00000063;
            8'd24: data = 32'h00000057;
            8'd25: data = 32'h0000004c;
            8'd26: data = 32'h00000058;
            8'd27: data = 32'h00000037;
            8'd28: data = 32'h00000063;
            8'd29: data = 32'h0000004d;
            8'd30: data = 32'h00000057;
            8'd31: data = 32'h00000061;
            8'd32: data = 32'h0000005f;
            8'd33: data = 32'h0000004d;
            8'd34: data = 32'h00000036;
            8'd35: data = 32'h00000063;
            8'd36: data = 32'h00000057;
            8'd37: data = 32'h00000063;
            8'd38: data = 32'h00000041;
            8'd39: data = 32'h0000004a;
            8'd40: data = 32'h00000061;
            8'd41: data = 32'h00000063;
            8'd42: data = 32'h00000057;
            8'd43: data = 32'h0000004d;
            8'd44: data = 32'h0000004d;
            8'd45: data = 32'h00000063;
            8'd46: data = 32'h0000004d;
            8'd47: data = 32'h00000056;
            8'd48: data = 32'h00000058;
            8'd49: data = 32'h00000062;
            8'd50: data = 32'h00000062;
            8'd51: data = 32'h0000004d;
            8'd52: data = 32'h00000062;
            8'd53: data = 32'h0000004d;
            8'd54: data = 32'h00000042;
            8'd55: data = 32'h00000060;
            8'd56: data = 32'h0000004d;
            8'd57: data = 32'h00000041;
            8'd58: data = 32'h0000004d;
            8'd59: data = 32'h00000063;
            8'd60: data = 32'h00000036;
            8'd61: data = 32'h0000004b;
            8'd62: data = 32'h00000060;
            8'd63: data = 32'h00000062;
            8'd64: data = 32'h00000055;
            8'd65: data = 32'h00000057;
            8'd66: data = 32'h0000005f;
            8'd67: data = 32'h00000058;
            8'd68: data = 32'h00000063;
            8'd69: data = 32'h00000063;
            8'd70: data = 32'h00000057;
            8'd71: data = 32'h0000002b;
            8'd72: data = 32'h0000005f;
            8'd73: data = 32'h00000037;
            8'd74: data = 32'h00000061;
            8'd75: data = 32'h0000004d;
            8'd76: data = 32'h0000002c;
            8'd77: data = 32'h00000057;
            8'd78: data = 32'h00000042;
            8'd79: data = 32'h00000058;
            8'd80: data = 32'h00000063;
            8'd81: data = 32'h0000004d;
            8'd82: data = 32'h00000058;
            8'd83: data = 32'h00000058;
            8'd84: data = 32'h00000057;
            8'd85: data = 32'h0000004d;
            8'd86: data = 32'h00000062;
            8'd87: data = 32'h00000042;
            8'd88: data = 32'h00000042;
            8'd89: data = 32'h00000063;
            8'd90: data = 32'h00000061;
            8'd91: data = 32'h0000002c;
            8'd92: data = 32'h00000063;
            8'd93: data = 32'h00000061;
            8'd94: data = 32'h00000063;
            8'd95: data = 32'h00000059;
            8'd96: data = 32'h00000042;
            8'd97: data = 32'h00000037;
            8'd98: data = 32'h00000058;
            8'd99: data = 32'h0000004b;
            8'd100: data = 32'h00000061;
            8'd101: data = 32'h0000004d;
            8'd102: data = 32'h00000063;
            8'd103: data = 32'h00000057;
            8'd104: data = 32'h0000004c;
            8'd105: data = 32'h00000063;
            8'd106: data = 32'h00000063;
            8'd107: data = 32'h00000058;
            8'd108: data = 32'h00000058;
            8'd109: data = 32'h00000063;
            8'd110: data = 32'h00000062;
            8'd111: data = 32'h00000058;
            8'd112: data = 32'h00000054;
            8'd113: data = 32'h00000056;
            8'd114: data = 32'h00000063;
            8'd115: data = 32'h00000063;
            8'd116: data = 32'h00000058;
            8'd117: data = 32'h00000042;
            8'd118: data = 32'h0000004d;
            8'd119: data = 32'h00000057;
            8'd120: data = 32'h00000042;
            8'd121: data = 32'h00000056;
            8'd122: data = 32'h00000063;
            8'd123: data = 32'h00000063;
            8'd124: data = 32'h0000004d;
            8'd125: data = 32'h0000004d;
            8'd126: data = 32'h00000057;
            8'd127: data = 32'h00000057;
            8'd128: data = 32'h00000060;
            8'd129: data = 32'h00000063;
            8'd130: data = 32'h00000061;
            8'd131: data = 32'h00000056;
            8'd132: data = 32'h00000063;
            8'd133: data = 32'h00000055;
            8'd134: data = 32'h00000037;
            8'd135: data = 32'h00000059;
            8'd136: data = 32'h00000058;
            8'd137: data = 32'h00000062;
            8'd138: data = 32'h0000004d;
            8'd139: data = 32'h00000056;
            8'd140: data = 32'h0000004d;
            8'd141: data = 32'h00000042;
            8'd142: data = 32'h00000061;
            8'd143: data = 32'h00000059;
            8'd144: data = 32'h00000056;
            8'd145: data = 32'h00000041;
            8'd146: data = 32'h00000041;
            8'd147: data = 32'h00000063;
            8'd148: data = 32'h00000063;
            8'd149: data = 32'h00000061;
            8'd150: data = 32'h00000058;
            8'd151: data = 32'h0000004a;
            8'd152: data = 32'h00000062;
            8'd153: data = 32'h00000063;
            8'd154: data = 32'h00000037;
            8'd155: data = 32'h00000057;
            8'd156: data = 32'h0000004d;
            8'd157: data = 32'h00000060;
            8'd158: data = 32'h0000002c;
            8'd159: data = 32'h00000058;
            8'd160: data = 32'h0000004d;
            8'd161: data = 32'h00000041;
            8'd162: data = 32'h00000060;
            8'd163: data = 32'h00000059;
            8'd164: data = 32'h00000057;
            8'd165: data = 32'h00000063;
            8'd166: data = 32'h00000057;
            8'd167: data = 32'h00000053;
            8'd168: data = 32'h00000056;
            8'd169: data = 32'h00000063;
            8'd170: data = 32'h00000057;
            8'd171: data = 32'h0000004c;
            8'd172: data = 32'h00000063;
            8'd173: data = 32'h00000063;
            8'd174: data = 32'h00000063;
            8'd175: data = 32'h00000059;
            8'd176: data = 32'h00000057;
            8'd177: data = 32'h00000062;
            8'd178: data = 32'h00000058;
            8'd179: data = 32'h0000004d;
            8'd180: data = 32'h00000063;
            8'd181: data = 32'h0000002c;
            8'd182: data = 32'h0000004d;
            8'd183: data = 32'h0000004d;
            8'd184: data = 32'h0000005f;
            8'd185: data = 32'h00000058;
            8'd186: data = 32'h0000004c;
            8'd187: data = 32'h0000004d;
            8'd188: data = 32'h0000004d;
            8'd189: data = 32'h0000004d;
            8'd190: data = 32'h0000004d;
            8'd191: data = 32'h00000063;
            8'd192: data = 32'h00000063;
            8'd193: data = 32'h0000004d;
            8'd194: data = 32'h00000056;
            8'd195: data = 32'h00000061;
            8'd196: data = 32'h00000057;
            8'd197: data = 32'h00000058;
            8'd198: data = 32'h00000037;
            8'd199: data = 32'h00000042;
            default: data = 32'b0;
        endcase
    end

endmodule
