localparam NUM_POINTS = 8;
