localparam NUM_NODES = 111;
localparam OUT_NODE = 0;
localparam YOU_NODE = 110;
