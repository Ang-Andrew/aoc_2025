localparam NUM_NODES = 1000;
localparam NUM_EDGES = 1000;
localparam K_LIMIT = 1000;
