// Day 5 ROM with match data
// Depth: 1000 entries (1000 IDs)
// Sum: 726

module rom_day5_data #(
    parameter WIDTH = 32,
    parameter DEPTH = 1000
) (
    input wire clk,
    input wire [9:0] addr,
    output reg [WIDTH-1:0] data
);

    reg [WIDTH-1:0] memory [0:DEPTH-1];

    initial begin
        // Initialize ROM with precomputed match data
        memory[   0] = 0;
        memory[   1] = 1;
        memory[   2] = 1;
        memory[   3] = 1;
        memory[   4] = 1;
        memory[   5] = 0;
        memory[   6] = 1;
        memory[   7] = 1;
        memory[   8] = 1;
        memory[   9] = 1;
        memory[  10] = 1;
        memory[  11] = 1;
        memory[  12] = 1;
        memory[  13] = 1;
        memory[  14] = 1;
        memory[  15] = 1;
        memory[  16] = 1;
        memory[  17] = 1;
        memory[  18] = 1;
        memory[  19] = 1;
        memory[  20] = 1;
        memory[  21] = 0;
        memory[  22] = 0;
        memory[  23] = 0;
        memory[  24] = 1;
        memory[  25] = 0;
        memory[  26] = 1;
        memory[  27] = 1;
        memory[  28] = 1;
        memory[  29] = 1;
        memory[  30] = 0;
        memory[  31] = 0;
        memory[  32] = 1;
        memory[  33] = 1;
        memory[  34] = 1;
        memory[  35] = 0;
        memory[  36] = 1;
        memory[  37] = 1;
        memory[  38] = 1;
        memory[  39] = 0;
        memory[  40] = 1;
        memory[  41] = 1;
        memory[  42] = 1;
        memory[  43] = 1;
        memory[  44] = 1;
        memory[  45] = 1;
        memory[  46] = 1;
        memory[  47] = 1;
        memory[  48] = 0;
        memory[  49] = 1;
        memory[  50] = 1;
        memory[  51] = 0;
        memory[  52] = 1;
        memory[  53] = 0;
        memory[  54] = 1;
        memory[  55] = 1;
        memory[  56] = 0;
        memory[  57] = 0;
        memory[  58] = 1;
        memory[  59] = 1;
        memory[  60] = 1;
        memory[  61] = 1;
        memory[  62] = 1;
        memory[  63] = 1;
        memory[  64] = 1;
        memory[  65] = 0;
        memory[  66] = 1;
        memory[  67] = 0;
        memory[  68] = 0;
        memory[  69] = 1;
        memory[  70] = 1;
        memory[  71] = 0;
        memory[  72] = 1;
        memory[  73] = 1;
        memory[  74] = 0;
        memory[  75] = 1;
        memory[  76] = 1;
        memory[  77] = 1;
        memory[  78] = 1;
        memory[  79] = 1;
        memory[  80] = 1;
        memory[  81] = 1;
        memory[  82] = 1;
        memory[  83] = 1;
        memory[  84] = 1;
        memory[  85] = 1;
        memory[  86] = 1;
        memory[  87] = 1;
        memory[  88] = 1;
        memory[  89] = 0;
        memory[  90] = 1;
        memory[  91] = 1;
        memory[  92] = 1;
        memory[  93] = 0;
        memory[  94] = 1;
        memory[  95] = 0;
        memory[  96] = 0;
        memory[  97] = 1;
        memory[  98] = 1;
        memory[  99] = 1;
        memory[ 100] = 1;
        memory[ 101] = 0;
        memory[ 102] = 0;
        memory[ 103] = 1;
        memory[ 104] = 1;
        memory[ 105] = 0;
        memory[ 106] = 0;
        memory[ 107] = 0;
        memory[ 108] = 1;
        memory[ 109] = 1;
        memory[ 110] = 1;
        memory[ 111] = 1;
        memory[ 112] = 1;
        memory[ 113] = 1;
        memory[ 114] = 0;
        memory[ 115] = 1;
        memory[ 116] = 1;
        memory[ 117] = 1;
        memory[ 118] = 0;
        memory[ 119] = 1;
        memory[ 120] = 0;
        memory[ 121] = 1;
        memory[ 122] = 1;
        memory[ 123] = 1;
        memory[ 124] = 1;
        memory[ 125] = 1;
        memory[ 126] = 1;
        memory[ 127] = 0;
        memory[ 128] = 1;
        memory[ 129] = 1;
        memory[ 130] = 1;
        memory[ 131] = 0;
        memory[ 132] = 1;
        memory[ 133] = 0;
        memory[ 134] = 0;
        memory[ 135] = 1;
        memory[ 136] = 1;
        memory[ 137] = 0;
        memory[ 138] = 1;
        memory[ 139] = 1;
        memory[ 140] = 1;
        memory[ 141] = 1;
        memory[ 142] = 1;
        memory[ 143] = 1;
        memory[ 144] = 0;
        memory[ 145] = 0;
        memory[ 146] = 0;
        memory[ 147] = 1;
        memory[ 148] = 0;
        memory[ 149] = 0;
        memory[ 150] = 1;
        memory[ 151] = 1;
        memory[ 152] = 0;
        memory[ 153] = 0;
        memory[ 154] = 1;
        memory[ 155] = 1;
        memory[ 156] = 1;
        memory[ 157] = 1;
        memory[ 158] = 1;
        memory[ 159] = 1;
        memory[ 160] = 1;
        memory[ 161] = 1;
        memory[ 162] = 0;
        memory[ 163] = 1;
        memory[ 164] = 1;
        memory[ 165] = 1;
        memory[ 166] = 0;
        memory[ 167] = 1;
        memory[ 168] = 1;
        memory[ 169] = 1;
        memory[ 170] = 1;
        memory[ 171] = 0;
        memory[ 172] = 1;
        memory[ 173] = 1;
        memory[ 174] = 1;
        memory[ 175] = 1;
        memory[ 176] = 1;
        memory[ 177] = 1;
        memory[ 178] = 0;
        memory[ 179] = 1;
        memory[ 180] = 1;
        memory[ 181] = 0;
        memory[ 182] = 1;
        memory[ 183] = 1;
        memory[ 184] = 1;
        memory[ 185] = 1;
        memory[ 186] = 0;
        memory[ 187] = 0;
        memory[ 188] = 0;
        memory[ 189] = 1;
        memory[ 190] = 1;
        memory[ 191] = 1;
        memory[ 192] = 1;
        memory[ 193] = 1;
        memory[ 194] = 1;
        memory[ 195] = 1;
        memory[ 196] = 1;
        memory[ 197] = 1;
        memory[ 198] = 1;
        memory[ 199] = 1;
        memory[ 200] = 1;
        memory[ 201] = 0;
        memory[ 202] = 1;
        memory[ 203] = 1;
        memory[ 204] = 1;
        memory[ 205] = 0;
        memory[ 206] = 1;
        memory[ 207] = 1;
        memory[ 208] = 1;
        memory[ 209] = 0;
        memory[ 210] = 1;
        memory[ 211] = 1;
        memory[ 212] = 1;
        memory[ 213] = 0;
        memory[ 214] = 1;
        memory[ 215] = 1;
        memory[ 216] = 1;
        memory[ 217] = 1;
        memory[ 218] = 0;
        memory[ 219] = 0;
        memory[ 220] = 1;
        memory[ 221] = 1;
        memory[ 222] = 1;
        memory[ 223] = 1;
        memory[ 224] = 1;
        memory[ 225] = 0;
        memory[ 226] = 1;
        memory[ 227] = 1;
        memory[ 228] = 1;
        memory[ 229] = 0;
        memory[ 230] = 1;
        memory[ 231] = 1;
        memory[ 232] = 1;
        memory[ 233] = 1;
        memory[ 234] = 0;
        memory[ 235] = 0;
        memory[ 236] = 1;
        memory[ 237] = 1;
        memory[ 238] = 1;
        memory[ 239] = 1;
        memory[ 240] = 0;
        memory[ 241] = 1;
        memory[ 242] = 0;
        memory[ 243] = 1;
        memory[ 244] = 1;
        memory[ 245] = 1;
        memory[ 246] = 1;
        memory[ 247] = 1;
        memory[ 248] = 1;
        memory[ 249] = 1;
        memory[ 250] = 0;
        memory[ 251] = 1;
        memory[ 252] = 1;
        memory[ 253] = 1;
        memory[ 254] = 1;
        memory[ 255] = 1;
        memory[ 256] = 0;
        memory[ 257] = 1;
        memory[ 258] = 1;
        memory[ 259] = 0;
        memory[ 260] = 1;
        memory[ 261] = 0;
        memory[ 262] = 1;
        memory[ 263] = 0;
        memory[ 264] = 1;
        memory[ 265] = 1;
        memory[ 266] = 1;
        memory[ 267] = 0;
        memory[ 268] = 1;
        memory[ 269] = 1;
        memory[ 270] = 1;
        memory[ 271] = 1;
        memory[ 272] = 1;
        memory[ 273] = 1;
        memory[ 274] = 1;
        memory[ 275] = 1;
        memory[ 276] = 0;
        memory[ 277] = 1;
        memory[ 278] = 0;
        memory[ 279] = 0;
        memory[ 280] = 0;
        memory[ 281] = 1;
        memory[ 282] = 1;
        memory[ 283] = 1;
        memory[ 284] = 1;
        memory[ 285] = 0;
        memory[ 286] = 1;
        memory[ 287] = 1;
        memory[ 288] = 1;
        memory[ 289] = 1;
        memory[ 290] = 0;
        memory[ 291] = 1;
        memory[ 292] = 0;
        memory[ 293] = 0;
        memory[ 294] = 1;
        memory[ 295] = 1;
        memory[ 296] = 1;
        memory[ 297] = 0;
        memory[ 298] = 1;
        memory[ 299] = 0;
        memory[ 300] = 1;
        memory[ 301] = 1;
        memory[ 302] = 1;
        memory[ 303] = 1;
        memory[ 304] = 1;
        memory[ 305] = 1;
        memory[ 306] = 1;
        memory[ 307] = 1;
        memory[ 308] = 1;
        memory[ 309] = 1;
        memory[ 310] = 1;
        memory[ 311] = 0;
        memory[ 312] = 1;
        memory[ 313] = 0;
        memory[ 314] = 1;
        memory[ 315] = 1;
        memory[ 316] = 0;
        memory[ 317] = 1;
        memory[ 318] = 1;
        memory[ 319] = 1;
        memory[ 320] = 1;
        memory[ 321] = 1;
        memory[ 322] = 1;
        memory[ 323] = 1;
        memory[ 324] = 1;
        memory[ 325] = 0;
        memory[ 326] = 1;
        memory[ 327] = 1;
        memory[ 328] = 0;
        memory[ 329] = 0;
        memory[ 330] = 1;
        memory[ 331] = 1;
        memory[ 332] = 0;
        memory[ 333] = 1;
        memory[ 334] = 1;
        memory[ 335] = 1;
        memory[ 336] = 1;
        memory[ 337] = 0;
        memory[ 338] = 0;
        memory[ 339] = 1;
        memory[ 340] = 1;
        memory[ 341] = 1;
        memory[ 342] = 1;
        memory[ 343] = 1;
        memory[ 344] = 1;
        memory[ 345] = 0;
        memory[ 346] = 1;
        memory[ 347] = 1;
        memory[ 348] = 0;
        memory[ 349] = 1;
        memory[ 350] = 1;
        memory[ 351] = 1;
        memory[ 352] = 1;
        memory[ 353] = 1;
        memory[ 354] = 1;
        memory[ 355] = 1;
        memory[ 356] = 1;
        memory[ 357] = 0;
        memory[ 358] = 1;
        memory[ 359] = 1;
        memory[ 360] = 1;
        memory[ 361] = 1;
        memory[ 362] = 0;
        memory[ 363] = 1;
        memory[ 364] = 1;
        memory[ 365] = 0;
        memory[ 366] = 1;
        memory[ 367] = 1;
        memory[ 368] = 0;
        memory[ 369] = 1;
        memory[ 370] = 1;
        memory[ 371] = 1;
        memory[ 372] = 1;
        memory[ 373] = 0;
        memory[ 374] = 1;
        memory[ 375] = 0;
        memory[ 376] = 1;
        memory[ 377] = 1;
        memory[ 378] = 1;
        memory[ 379] = 0;
        memory[ 380] = 1;
        memory[ 381] = 0;
        memory[ 382] = 1;
        memory[ 383] = 0;
        memory[ 384] = 1;
        memory[ 385] = 0;
        memory[ 386] = 1;
        memory[ 387] = 1;
        memory[ 388] = 0;
        memory[ 389] = 0;
        memory[ 390] = 1;
        memory[ 391] = 0;
        memory[ 392] = 1;
        memory[ 393] = 1;
        memory[ 394] = 1;
        memory[ 395] = 0;
        memory[ 396] = 0;
        memory[ 397] = 1;
        memory[ 398] = 1;
        memory[ 399] = 1;
        memory[ 400] = 0;
        memory[ 401] = 1;
        memory[ 402] = 0;
        memory[ 403] = 0;
        memory[ 404] = 0;
        memory[ 405] = 1;
        memory[ 406] = 0;
        memory[ 407] = 0;
        memory[ 408] = 1;
        memory[ 409] = 1;
        memory[ 410] = 1;
        memory[ 411] = 1;
        memory[ 412] = 1;
        memory[ 413] = 1;
        memory[ 414] = 1;
        memory[ 415] = 1;
        memory[ 416] = 1;
        memory[ 417] = 0;
        memory[ 418] = 1;
        memory[ 419] = 1;
        memory[ 420] = 1;
        memory[ 421] = 0;
        memory[ 422] = 1;
        memory[ 423] = 1;
        memory[ 424] = 1;
        memory[ 425] = 1;
        memory[ 426] = 1;
        memory[ 427] = 1;
        memory[ 428] = 1;
        memory[ 429] = 0;
        memory[ 430] = 1;
        memory[ 431] = 1;
        memory[ 432] = 1;
        memory[ 433] = 0;
        memory[ 434] = 1;
        memory[ 435] = 1;
        memory[ 436] = 0;
        memory[ 437] = 1;
        memory[ 438] = 1;
        memory[ 439] = 1;
        memory[ 440] = 1;
        memory[ 441] = 1;
        memory[ 442] = 1;
        memory[ 443] = 1;
        memory[ 444] = 1;
        memory[ 445] = 1;
        memory[ 446] = 1;
        memory[ 447] = 1;
        memory[ 448] = 1;
        memory[ 449] = 0;
        memory[ 450] = 1;
        memory[ 451] = 0;
        memory[ 452] = 1;
        memory[ 453] = 0;
        memory[ 454] = 1;
        memory[ 455] = 1;
        memory[ 456] = 1;
        memory[ 457] = 1;
        memory[ 458] = 1;
        memory[ 459] = 0;
        memory[ 460] = 1;
        memory[ 461] = 1;
        memory[ 462] = 1;
        memory[ 463] = 1;
        memory[ 464] = 1;
        memory[ 465] = 1;
        memory[ 466] = 1;
        memory[ 467] = 1;
        memory[ 468] = 0;
        memory[ 469] = 0;
        memory[ 470] = 1;
        memory[ 471] = 1;
        memory[ 472] = 1;
        memory[ 473] = 1;
        memory[ 474] = 1;
        memory[ 475] = 0;
        memory[ 476] = 1;
        memory[ 477] = 1;
        memory[ 478] = 0;
        memory[ 479] = 1;
        memory[ 480] = 1;
        memory[ 481] = 1;
        memory[ 482] = 1;
        memory[ 483] = 1;
        memory[ 484] = 0;
        memory[ 485] = 1;
        memory[ 486] = 0;
        memory[ 487] = 0;
        memory[ 488] = 0;
        memory[ 489] = 1;
        memory[ 490] = 0;
        memory[ 491] = 0;
        memory[ 492] = 1;
        memory[ 493] = 1;
        memory[ 494] = 1;
        memory[ 495] = 1;
        memory[ 496] = 1;
        memory[ 497] = 1;
        memory[ 498] = 1;
        memory[ 499] = 1;
        memory[ 500] = 0;
        memory[ 501] = 1;
        memory[ 502] = 1;
        memory[ 503] = 1;
        memory[ 504] = 1;
        memory[ 505] = 1;
        memory[ 506] = 0;
        memory[ 507] = 1;
        memory[ 508] = 1;
        memory[ 509] = 1;
        memory[ 510] = 1;
        memory[ 511] = 1;
        memory[ 512] = 0;
        memory[ 513] = 1;
        memory[ 514] = 1;
        memory[ 515] = 0;
        memory[ 516] = 1;
        memory[ 517] = 1;
        memory[ 518] = 0;
        memory[ 519] = 1;
        memory[ 520] = 1;
        memory[ 521] = 0;
        memory[ 522] = 1;
        memory[ 523] = 1;
        memory[ 524] = 1;
        memory[ 525] = 1;
        memory[ 526] = 1;
        memory[ 527] = 0;
        memory[ 528] = 0;
        memory[ 529] = 1;
        memory[ 530] = 0;
        memory[ 531] = 1;
        memory[ 532] = 1;
        memory[ 533] = 1;
        memory[ 534] = 1;
        memory[ 535] = 1;
        memory[ 536] = 0;
        memory[ 537] = 1;
        memory[ 538] = 0;
        memory[ 539] = 1;
        memory[ 540] = 1;
        memory[ 541] = 0;
        memory[ 542] = 1;
        memory[ 543] = 0;
        memory[ 544] = 1;
        memory[ 545] = 1;
        memory[ 546] = 1;
        memory[ 547] = 0;
        memory[ 548] = 1;
        memory[ 549] = 1;
        memory[ 550] = 1;
        memory[ 551] = 0;
        memory[ 552] = 1;
        memory[ 553] = 1;
        memory[ 554] = 0;
        memory[ 555] = 0;
        memory[ 556] = 0;
        memory[ 557] = 1;
        memory[ 558] = 1;
        memory[ 559] = 1;
        memory[ 560] = 1;
        memory[ 561] = 0;
        memory[ 562] = 0;
        memory[ 563] = 0;
        memory[ 564] = 1;
        memory[ 565] = 1;
        memory[ 566] = 1;
        memory[ 567] = 1;
        memory[ 568] = 1;
        memory[ 569] = 1;
        memory[ 570] = 1;
        memory[ 571] = 0;
        memory[ 572] = 0;
        memory[ 573] = 1;
        memory[ 574] = 1;
        memory[ 575] = 0;
        memory[ 576] = 1;
        memory[ 577] = 1;
        memory[ 578] = 1;
        memory[ 579] = 1;
        memory[ 580] = 1;
        memory[ 581] = 1;
        memory[ 582] = 1;
        memory[ 583] = 1;
        memory[ 584] = 0;
        memory[ 585] = 0;
        memory[ 586] = 1;
        memory[ 587] = 1;
        memory[ 588] = 0;
        memory[ 589] = 1;
        memory[ 590] = 1;
        memory[ 591] = 1;
        memory[ 592] = 1;
        memory[ 593] = 0;
        memory[ 594] = 1;
        memory[ 595] = 1;
        memory[ 596] = 1;
        memory[ 597] = 1;
        memory[ 598] = 1;
        memory[ 599] = 1;
        memory[ 600] = 1;
        memory[ 601] = 0;
        memory[ 602] = 1;
        memory[ 603] = 0;
        memory[ 604] = 0;
        memory[ 605] = 0;
        memory[ 606] = 1;
        memory[ 607] = 1;
        memory[ 608] = 1;
        memory[ 609] = 1;
        memory[ 610] = 1;
        memory[ 611] = 1;
        memory[ 612] = 1;
        memory[ 613] = 1;
        memory[ 614] = 0;
        memory[ 615] = 0;
        memory[ 616] = 1;
        memory[ 617] = 0;
        memory[ 618] = 0;
        memory[ 619] = 1;
        memory[ 620] = 1;
        memory[ 621] = 1;
        memory[ 622] = 0;
        memory[ 623] = 0;
        memory[ 624] = 0;
        memory[ 625] = 1;
        memory[ 626] = 1;
        memory[ 627] = 1;
        memory[ 628] = 0;
        memory[ 629] = 1;
        memory[ 630] = 1;
        memory[ 631] = 0;
        memory[ 632] = 1;
        memory[ 633] = 1;
        memory[ 634] = 1;
        memory[ 635] = 1;
        memory[ 636] = 1;
        memory[ 637] = 1;
        memory[ 638] = 0;
        memory[ 639] = 1;
        memory[ 640] = 0;
        memory[ 641] = 0;
        memory[ 642] = 1;
        memory[ 643] = 0;
        memory[ 644] = 1;
        memory[ 645] = 1;
        memory[ 646] = 1;
        memory[ 647] = 0;
        memory[ 648] = 0;
        memory[ 649] = 0;
        memory[ 650] = 0;
        memory[ 651] = 1;
        memory[ 652] = 1;
        memory[ 653] = 1;
        memory[ 654] = 1;
        memory[ 655] = 1;
        memory[ 656] = 0;
        memory[ 657] = 1;
        memory[ 658] = 1;
        memory[ 659] = 0;
        memory[ 660] = 1;
        memory[ 661] = 1;
        memory[ 662] = 1;
        memory[ 663] = 0;
        memory[ 664] = 1;
        memory[ 665] = 1;
        memory[ 666] = 1;
        memory[ 667] = 1;
        memory[ 668] = 0;
        memory[ 669] = 1;
        memory[ 670] = 1;
        memory[ 671] = 1;
        memory[ 672] = 1;
        memory[ 673] = 1;
        memory[ 674] = 0;
        memory[ 675] = 1;
        memory[ 676] = 1;
        memory[ 677] = 1;
        memory[ 678] = 1;
        memory[ 679] = 0;
        memory[ 680] = 1;
        memory[ 681] = 0;
        memory[ 682] = 0;
        memory[ 683] = 1;
        memory[ 684] = 0;
        memory[ 685] = 0;
        memory[ 686] = 1;
        memory[ 687] = 0;
        memory[ 688] = 1;
        memory[ 689] = 1;
        memory[ 690] = 1;
        memory[ 691] = 1;
        memory[ 692] = 1;
        memory[ 693] = 1;
        memory[ 694] = 1;
        memory[ 695] = 1;
        memory[ 696] = 1;
        memory[ 697] = 0;
        memory[ 698] = 1;
        memory[ 699] = 1;
        memory[ 700] = 1;
        memory[ 701] = 0;
        memory[ 702] = 1;
        memory[ 703] = 0;
        memory[ 704] = 1;
        memory[ 705] = 0;
        memory[ 706] = 0;
        memory[ 707] = 1;
        memory[ 708] = 0;
        memory[ 709] = 1;
        memory[ 710] = 1;
        memory[ 711] = 0;
        memory[ 712] = 1;
        memory[ 713] = 1;
        memory[ 714] = 1;
        memory[ 715] = 1;
        memory[ 716] = 0;
        memory[ 717] = 0;
        memory[ 718] = 1;
        memory[ 719] = 1;
        memory[ 720] = 1;
        memory[ 721] = 1;
        memory[ 722] = 1;
        memory[ 723] = 1;
        memory[ 724] = 0;
        memory[ 725] = 0;
        memory[ 726] = 1;
        memory[ 727] = 1;
        memory[ 728] = 1;
        memory[ 729] = 1;
        memory[ 730] = 0;
        memory[ 731] = 1;
        memory[ 732] = 1;
        memory[ 733] = 1;
        memory[ 734] = 0;
        memory[ 735] = 1;
        memory[ 736] = 1;
        memory[ 737] = 0;
        memory[ 738] = 1;
        memory[ 739] = 1;
        memory[ 740] = 1;
        memory[ 741] = 1;
        memory[ 742] = 0;
        memory[ 743] = 1;
        memory[ 744] = 1;
        memory[ 745] = 1;
        memory[ 746] = 1;
        memory[ 747] = 1;
        memory[ 748] = 0;
        memory[ 749] = 0;
        memory[ 750] = 0;
        memory[ 751] = 1;
        memory[ 752] = 1;
        memory[ 753] = 1;
        memory[ 754] = 1;
        memory[ 755] = 1;
        memory[ 756] = 1;
        memory[ 757] = 0;
        memory[ 758] = 1;
        memory[ 759] = 1;
        memory[ 760] = 1;
        memory[ 761] = 1;
        memory[ 762] = 1;
        memory[ 763] = 1;
        memory[ 764] = 1;
        memory[ 765] = 1;
        memory[ 766] = 1;
        memory[ 767] = 1;
        memory[ 768] = 1;
        memory[ 769] = 1;
        memory[ 770] = 1;
        memory[ 771] = 1;
        memory[ 772] = 1;
        memory[ 773] = 1;
        memory[ 774] = 0;
        memory[ 775] = 1;
        memory[ 776] = 0;
        memory[ 777] = 1;
        memory[ 778] = 1;
        memory[ 779] = 1;
        memory[ 780] = 0;
        memory[ 781] = 1;
        memory[ 782] = 1;
        memory[ 783] = 0;
        memory[ 784] = 1;
        memory[ 785] = 1;
        memory[ 786] = 0;
        memory[ 787] = 1;
        memory[ 788] = 1;
        memory[ 789] = 1;
        memory[ 790] = 1;
        memory[ 791] = 1;
        memory[ 792] = 0;
        memory[ 793] = 1;
        memory[ 794] = 0;
        memory[ 795] = 1;
        memory[ 796] = 0;
        memory[ 797] = 1;
        memory[ 798] = 1;
        memory[ 799] = 1;
        memory[ 800] = 0;
        memory[ 801] = 0;
        memory[ 802] = 1;
        memory[ 803] = 1;
        memory[ 804] = 1;
        memory[ 805] = 1;
        memory[ 806] = 0;
        memory[ 807] = 1;
        memory[ 808] = 1;
        memory[ 809] = 1;
        memory[ 810] = 1;
        memory[ 811] = 1;
        memory[ 812] = 1;
        memory[ 813] = 1;
        memory[ 814] = 0;
        memory[ 815] = 0;
        memory[ 816] = 1;
        memory[ 817] = 0;
        memory[ 818] = 1;
        memory[ 819] = 1;
        memory[ 820] = 0;
        memory[ 821] = 1;
        memory[ 822] = 1;
        memory[ 823] = 1;
        memory[ 824] = 0;
        memory[ 825] = 0;
        memory[ 826] = 1;
        memory[ 827] = 1;
        memory[ 828] = 0;
        memory[ 829] = 0;
        memory[ 830] = 1;
        memory[ 831] = 1;
        memory[ 832] = 1;
        memory[ 833] = 1;
        memory[ 834] = 1;
        memory[ 835] = 0;
        memory[ 836] = 0;
        memory[ 837] = 1;
        memory[ 838] = 0;
        memory[ 839] = 1;
        memory[ 840] = 1;
        memory[ 841] = 1;
        memory[ 842] = 1;
        memory[ 843] = 1;
        memory[ 844] = 0;
        memory[ 845] = 0;
        memory[ 846] = 1;
        memory[ 847] = 1;
        memory[ 848] = 1;
        memory[ 849] = 1;
        memory[ 850] = 1;
        memory[ 851] = 1;
        memory[ 852] = 1;
        memory[ 853] = 1;
        memory[ 854] = 1;
        memory[ 855] = 1;
        memory[ 856] = 1;
        memory[ 857] = 1;
        memory[ 858] = 0;
        memory[ 859] = 1;
        memory[ 860] = 1;
        memory[ 861] = 1;
        memory[ 862] = 1;
        memory[ 863] = 1;
        memory[ 864] = 1;
        memory[ 865] = 1;
        memory[ 866] = 0;
        memory[ 867] = 0;
        memory[ 868] = 0;
        memory[ 869] = 0;
        memory[ 870] = 1;
        memory[ 871] = 1;
        memory[ 872] = 1;
        memory[ 873] = 1;
        memory[ 874] = 1;
        memory[ 875] = 0;
        memory[ 876] = 1;
        memory[ 877] = 1;
        memory[ 878] = 0;
        memory[ 879] = 1;
        memory[ 880] = 1;
        memory[ 881] = 1;
        memory[ 882] = 0;
        memory[ 883] = 1;
        memory[ 884] = 1;
        memory[ 885] = 1;
        memory[ 886] = 1;
        memory[ 887] = 1;
        memory[ 888] = 1;
        memory[ 889] = 1;
        memory[ 890] = 0;
        memory[ 891] = 1;
        memory[ 892] = 1;
        memory[ 893] = 1;
        memory[ 894] = 1;
        memory[ 895] = 0;
        memory[ 896] = 1;
        memory[ 897] = 1;
        memory[ 898] = 1;
        memory[ 899] = 1;
        memory[ 900] = 1;
        memory[ 901] = 0;
        memory[ 902] = 1;
        memory[ 903] = 1;
        memory[ 904] = 0;
        memory[ 905] = 1;
        memory[ 906] = 0;
        memory[ 907] = 1;
        memory[ 908] = 1;
        memory[ 909] = 0;
        memory[ 910] = 1;
        memory[ 911] = 1;
        memory[ 912] = 0;
        memory[ 913] = 1;
        memory[ 914] = 1;
        memory[ 915] = 1;
        memory[ 916] = 1;
        memory[ 917] = 0;
        memory[ 918] = 1;
        memory[ 919] = 0;
        memory[ 920] = 1;
        memory[ 921] = 1;
        memory[ 922] = 0;
        memory[ 923] = 1;
        memory[ 924] = 1;
        memory[ 925] = 0;
        memory[ 926] = 1;
        memory[ 927] = 0;
        memory[ 928] = 1;
        memory[ 929] = 1;
        memory[ 930] = 1;
        memory[ 931] = 1;
        memory[ 932] = 0;
        memory[ 933] = 1;
        memory[ 934] = 1;
        memory[ 935] = 0;
        memory[ 936] = 1;
        memory[ 937] = 0;
        memory[ 938] = 1;
        memory[ 939] = 1;
        memory[ 940] = 1;
        memory[ 941] = 0;
        memory[ 942] = 1;
        memory[ 943] = 0;
        memory[ 944] = 1;
        memory[ 945] = 1;
        memory[ 946] = 0;
        memory[ 947] = 1;
        memory[ 948] = 1;
        memory[ 949] = 1;
        memory[ 950] = 0;
        memory[ 951] = 1;
        memory[ 952] = 1;
        memory[ 953] = 0;
        memory[ 954] = 1;
        memory[ 955] = 1;
        memory[ 956] = 1;
        memory[ 957] = 1;
        memory[ 958] = 0;
        memory[ 959] = 1;
        memory[ 960] = 1;
        memory[ 961] = 1;
        memory[ 962] = 1;
        memory[ 963] = 1;
        memory[ 964] = 1;
        memory[ 965] = 1;
        memory[ 966] = 0;
        memory[ 967] = 1;
        memory[ 968] = 0;
        memory[ 969] = 1;
        memory[ 970] = 1;
        memory[ 971] = 1;
        memory[ 972] = 0;
        memory[ 973] = 1;
        memory[ 974] = 1;
        memory[ 975] = 0;
        memory[ 976] = 0;
        memory[ 977] = 1;
        memory[ 978] = 1;
        memory[ 979] = 1;
        memory[ 980] = 1;
        memory[ 981] = 1;
        memory[ 982] = 0;
        memory[ 983] = 0;
        memory[ 984] = 1;
        memory[ 985] = 0;
        memory[ 986] = 1;
        memory[ 987] = 0;
        memory[ 988] = 1;
        memory[ 989] = 1;
        memory[ 990] = 1;
        memory[ 991] = 1;
        memory[ 992] = 1;
        memory[ 993] = 1;
        memory[ 994] = 1;
        memory[ 995] = 1;
        memory[ 996] = 0;
        memory[ 997] = 0;
        memory[ 998] = 1;
        memory[ 999] = 1;
    end

    always @(posedge clk) begin
        data <= memory[addr];
    end

endmodule
