localparam WIDTH = 141;
localparam HEIGHT = 142;
localparam MEM_SIZE = 20022;
