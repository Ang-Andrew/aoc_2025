localparam WIDTH = 15;
localparam HEIGHT = 16;
localparam MEM_SIZE = 240;
