localparam N = 1000;
localparam K = 10;
