// Day 4 ROM with hardcoded neighbor count data
// Depth: 12224 entries
// Sum: 1424

module rom_day4_hardcoded #(
    parameter WIDTH = 32,
    parameter DEPTH = 12224
) (
    input wire clk,
    input wire [13:0] addr,
    output reg [WIDTH-1:0] data
);

    reg [WIDTH-1:0] memory [0:DEPTH-1];

    initial begin
        // Initialize ROM with precomputed neighbor counts
        memory[    0] = 1;
        memory[    1] = 1;
        memory[    2] = 1;
        memory[    3] = 1;
        memory[    4] = 0;
        memory[    5] = 1;
        memory[    6] = 1;
        memory[    7] = 0;
        memory[    8] = 0;
        memory[    9] = 0;
        memory[   10] = 0;
        memory[   11] = 1;
        memory[   12] = 1;
        memory[   13] = 0;
        memory[   14] = 0;
        memory[   15] = 0;
        memory[   16] = 1;
        memory[   17] = 1;
        memory[   18] = 1;
        memory[   19] = 0;
        memory[   20] = 0;
        memory[   21] = 0;
        memory[   22] = 0;
        memory[   23] = 0;
        memory[   24] = 1;
        memory[   25] = 1;
        memory[   26] = 1;
        memory[   27] = 1;
        memory[   28] = 1;
        memory[   29] = 1;
        memory[   30] = 1;
        memory[   31] = 1;
        memory[   32] = 1;
        memory[   33] = 1;
        memory[   34] = 1;
        memory[   35] = 1;
        memory[   36] = 1;
        memory[   37] = 1;
        memory[   38] = 1;
        memory[   39] = 1;
        memory[   40] = 1;
        memory[   41] = 1;
        memory[   42] = 1;
        memory[   43] = 0;
        memory[   44] = 1;
        memory[   45] = 1;
        memory[   46] = 0;
        memory[   47] = 0;
        memory[   48] = 0;
        memory[   49] = 1;
        memory[   50] = 1;
        memory[   51] = 0;
        memory[   52] = 0;
        memory[   53] = 1;
        memory[   54] = 1;
        memory[   55] = 1;
        memory[   56] = 1;
        memory[   57] = 1;
        memory[   58] = 1;
        memory[   59] = 1;
        memory[   60] = 1;
        memory[   61] = 0;
        memory[   62] = 0;
        memory[   63] = 1;
        memory[   64] = 1;
        memory[   65] = 0;
        memory[   66] = 0;
        memory[   67] = 0;
        memory[   68] = 1;
        memory[   69] = 1;
        memory[   70] = 1;
        memory[   71] = 1;
        memory[   72] = 1;
        memory[   73] = 0;
        memory[   74] = 0;
        memory[   75] = 0;
        memory[   76] = 0;
        memory[   77] = 1;
        memory[   78] = 0;
        memory[   79] = 0;
        memory[   80] = 1;
        memory[   81] = 1;
        memory[   82] = 1;
        memory[   83] = 1;
        memory[   84] = 1;
        memory[   85] = 1;
        memory[   86] = 1;
        memory[   87] = 0;
        memory[   88] = 0;
        memory[   89] = 0;
        memory[   90] = 0;
        memory[   91] = 0;
        memory[   92] = 0;
        memory[   93] = 0;
        memory[   94] = 0;
        memory[   95] = 0;
        memory[   96] = 0;
        memory[   97] = 0;
        memory[   98] = 0;
        memory[   99] = 0;
        memory[  100] = 0;
        memory[  101] = 1;
        memory[  102] = 0;
        memory[  103] = 1;
        memory[  104] = 0;
        memory[  105] = 0;
        memory[  106] = 0;
        memory[  107] = 0;
        memory[  108] = 0;
        memory[  109] = 0;
        memory[  110] = 0;
        memory[  111] = 0;
        memory[  112] = 0;
        memory[  113] = 0;
        memory[  114] = 0;
        memory[  115] = 0;
        memory[  116] = 0;
        memory[  117] = 1;
        memory[  118] = 0;
        memory[  119] = 0;
        memory[  120] = 0;
        memory[  121] = 0;
        memory[  122] = 0;
        memory[  123] = 1;
        memory[  124] = 0;
        memory[  125] = 0;
        memory[  126] = 0;
        memory[  127] = 0;
        memory[  128] = 0;
        memory[  129] = 0;
        memory[  130] = 0;
        memory[  131] = 0;
        memory[  132] = 1;
        memory[  133] = 0;
        memory[  134] = 0;
        memory[  135] = 0;
        memory[  136] = 0;
        memory[  137] = 0;
        memory[  138] = 0;
        memory[  139] = 1;
        memory[  140] = 0;
        memory[  141] = 0;
        memory[  142] = 0;
        memory[  143] = 0;
        memory[  144] = 0;
        memory[  145] = 0;
        memory[  146] = 0;
        memory[  147] = 0;
        memory[  148] = 0;
        memory[  149] = 0;
        memory[  150] = 0;
        memory[  151] = 0;
        memory[  152] = 0;
        memory[  153] = 0;
        memory[  154] = 0;
        memory[  155] = 1;
        memory[  156] = 0;
        memory[  157] = 0;
        memory[  158] = 0;
        memory[  159] = 0;
        memory[  160] = 0;
        memory[  161] = 0;
        memory[  162] = 0;
        memory[  163] = 0;
        memory[  164] = 0;
        memory[  165] = 0;
        memory[  166] = 0;
        memory[  167] = 1;
        memory[  168] = 1;
        memory[  169] = 0;
        memory[  170] = 0;
        memory[  171] = 0;
        memory[  172] = 0;
        memory[  173] = 1;
        memory[  174] = 0;
        memory[  175] = 0;
        memory[  176] = 0;
        memory[  177] = 1;
        memory[  178] = 0;
        memory[  179] = 0;
        memory[  180] = 0;
        memory[  181] = 0;
        memory[  182] = 0;
        memory[  183] = 0;
        memory[  184] = 0;
        memory[  185] = 0;
        memory[  186] = 0;
        memory[  187] = 0;
        memory[  188] = 0;
        memory[  189] = 0;
        memory[  190] = 0;
        memory[  191] = 0;
        memory[  192] = 0;
        memory[  193] = 0;
        memory[  194] = 0;
        memory[  195] = 0;
        memory[  196] = 0;
        memory[  197] = 0;
        memory[  198] = 0;
        memory[  199] = 0;
        memory[  200] = 0;
        memory[  201] = 0;
        memory[  202] = 0;
        memory[  203] = 1;
        memory[  204] = 1;
        memory[  205] = 0;
        memory[  206] = 0;
        memory[  207] = 1;
        memory[  208] = 0;
        memory[  209] = 0;
        memory[  210] = 0;
        memory[  211] = 0;
        memory[  212] = 0;
        memory[  213] = 0;
        memory[  214] = 0;
        memory[  215] = 0;
        memory[  216] = 0;
        memory[  217] = 0;
        memory[  218] = 0;
        memory[  219] = 0;
        memory[  220] = 0;
        memory[  221] = 0;
        memory[  222] = 0;
        memory[  223] = 0;
        memory[  224] = 0;
        memory[  225] = 0;
        memory[  226] = 0;
        memory[  227] = 0;
        memory[  228] = 0;
        memory[  229] = 0;
        memory[  230] = 0;
        memory[  231] = 0;
        memory[  232] = 0;
        memory[  233] = 0;
        memory[  234] = 0;
        memory[  235] = 0;
        memory[  236] = 0;
        memory[  237] = 0;
        memory[  238] = 0;
        memory[  239] = 1;
        memory[  240] = 0;
        memory[  241] = 0;
        memory[  242] = 0;
        memory[  243] = 0;
        memory[  244] = 0;
        memory[  245] = 0;
        memory[  246] = 0;
        memory[  247] = 0;
        memory[  248] = 0;
        memory[  249] = 1;
        memory[  250] = 0;
        memory[  251] = 0;
        memory[  252] = 0;
        memory[  253] = 0;
        memory[  254] = 0;
        memory[  255] = 0;
        memory[  256] = 0;
        memory[  257] = 0;
        memory[  258] = 0;
        memory[  259] = 0;
        memory[  260] = 0;
        memory[  261] = 0;
        memory[  262] = 0;
        memory[  263] = 0;
        memory[  264] = 0;
        memory[  265] = 0;
        memory[  266] = 0;
        memory[  267] = 0;
        memory[  268] = 1;
        memory[  269] = 0;
        memory[  270] = 0;
        memory[  271] = 0;
        memory[  272] = 1;
        memory[  273] = 1;
        memory[  274] = 0;
        memory[  275] = 0;
        memory[  276] = 0;
        memory[  277] = 0;
        memory[  278] = 0;
        memory[  279] = 0;
        memory[  280] = 0;
        memory[  281] = 0;
        memory[  282] = 0;
        memory[  283] = 0;
        memory[  284] = 0;
        memory[  285] = 0;
        memory[  286] = 0;
        memory[  287] = 0;
        memory[  288] = 0;
        memory[  289] = 0;
        memory[  290] = 0;
        memory[  291] = 0;
        memory[  292] = 0;
        memory[  293] = 0;
        memory[  294] = 0;
        memory[  295] = 0;
        memory[  296] = 0;
        memory[  297] = 0;
        memory[  298] = 0;
        memory[  299] = 0;
        memory[  300] = 0;
        memory[  301] = 0;
        memory[  302] = 0;
        memory[  303] = 0;
        memory[  304] = 0;
        memory[  305] = 0;
        memory[  306] = 0;
        memory[  307] = 0;
        memory[  308] = 0;
        memory[  309] = 0;
        memory[  310] = 0;
        memory[  311] = 0;
        memory[  312] = 0;
        memory[  313] = 0;
        memory[  314] = 0;
        memory[  315] = 0;
        memory[  316] = 1;
        memory[  317] = 0;
        memory[  318] = 0;
        memory[  319] = 0;
        memory[  320] = 0;
        memory[  321] = 0;
        memory[  322] = 0;
        memory[  323] = 0;
        memory[  324] = 0;
        memory[  325] = 0;
        memory[  326] = 0;
        memory[  327] = 0;
        memory[  328] = 0;
        memory[  329] = 0;
        memory[  330] = 0;
        memory[  331] = 0;
        memory[  332] = 0;
        memory[  333] = 0;
        memory[  334] = 1;
        memory[  335] = 0;
        memory[  336] = 0;
        memory[  337] = 0;
        memory[  338] = 1;
        memory[  339] = 0;
        memory[  340] = 0;
        memory[  341] = 0;
        memory[  342] = 0;
        memory[  343] = 0;
        memory[  344] = 0;
        memory[  345] = 0;
        memory[  346] = 1;
        memory[  347] = 1;
        memory[  348] = 0;
        memory[  349] = 0;
        memory[  350] = 0;
        memory[  351] = 0;
        memory[  352] = 0;
        memory[  353] = 0;
        memory[  354] = 1;
        memory[  355] = 1;
        memory[  356] = 0;
        memory[  357] = 0;
        memory[  358] = 0;
        memory[  359] = 0;
        memory[  360] = 0;
        memory[  361] = 1;
        memory[  362] = 1;
        memory[  363] = 0;
        memory[  364] = 0;
        memory[  365] = 0;
        memory[  366] = 0;
        memory[  367] = 0;
        memory[  368] = 0;
        memory[  369] = 0;
        memory[  370] = 0;
        memory[  371] = 0;
        memory[  372] = 0;
        memory[  373] = 0;
        memory[  374] = 0;
        memory[  375] = 0;
        memory[  376] = 0;
        memory[  377] = 0;
        memory[  378] = 0;
        memory[  379] = 0;
        memory[  380] = 0;
        memory[  381] = 0;
        memory[  382] = 0;
        memory[  383] = 0;
        memory[  384] = 0;
        memory[  385] = 0;
        memory[  386] = 0;
        memory[  387] = 0;
        memory[  388] = 0;
        memory[  389] = 0;
        memory[  390] = 0;
        memory[  391] = 0;
        memory[  392] = 0;
        memory[  393] = 0;
        memory[  394] = 0;
        memory[  395] = 0;
        memory[  396] = 0;
        memory[  397] = 0;
        memory[  398] = 1;
        memory[  399] = 0;
        memory[  400] = 0;
        memory[  401] = 0;
        memory[  402] = 0;
        memory[  403] = 0;
        memory[  404] = 0;
        memory[  405] = 0;
        memory[  406] = 0;
        memory[  407] = 0;
        memory[  408] = 0;
        memory[  409] = 0;
        memory[  410] = 0;
        memory[  411] = 0;
        memory[  412] = 1;
        memory[  413] = 0;
        memory[  414] = 0;
        memory[  415] = 0;
        memory[  416] = 1;
        memory[  417] = 0;
        memory[  418] = 0;
        memory[  419] = 0;
        memory[  420] = 0;
        memory[  421] = 0;
        memory[  422] = 0;
        memory[  423] = 0;
        memory[  424] = 0;
        memory[  425] = 0;
        memory[  426] = 0;
        memory[  427] = 0;
        memory[  428] = 0;
        memory[  429] = 0;
        memory[  430] = 0;
        memory[  431] = 0;
        memory[  432] = 0;
        memory[  433] = 0;
        memory[  434] = 0;
        memory[  435] = 0;
        memory[  436] = 0;
        memory[  437] = 0;
        memory[  438] = 0;
        memory[  439] = 0;
        memory[  440] = 0;
        memory[  441] = 0;
        memory[  442] = 0;
        memory[  443] = 0;
        memory[  444] = 0;
        memory[  445] = 0;
        memory[  446] = 0;
        memory[  447] = 0;
        memory[  448] = 0;
        memory[  449] = 0;
        memory[  450] = 1;
        memory[  451] = 0;
        memory[  452] = 0;
        memory[  453] = 1;
        memory[  454] = 0;
        memory[  455] = 0;
        memory[  456] = 0;
        memory[  457] = 0;
        memory[  458] = 0;
        memory[  459] = 0;
        memory[  460] = 0;
        memory[  461] = 0;
        memory[  462] = 0;
        memory[  463] = 0;
        memory[  464] = 0;
        memory[  465] = 0;
        memory[  466] = 0;
        memory[  467] = 0;
        memory[  468] = 0;
        memory[  469] = 0;
        memory[  470] = 0;
        memory[  471] = 0;
        memory[  472] = 0;
        memory[  473] = 0;
        memory[  474] = 0;
        memory[  475] = 0;
        memory[  476] = 0;
        memory[  477] = 0;
        memory[  478] = 0;
        memory[  479] = 0;
        memory[  480] = 0;
        memory[  481] = 1;
        memory[  482] = 1;
        memory[  483] = 0;
        memory[  484] = 0;
        memory[  485] = 0;
        memory[  486] = 0;
        memory[  487] = 0;
        memory[  488] = 0;
        memory[  489] = 0;
        memory[  490] = 0;
        memory[  491] = 0;
        memory[  492] = 0;
        memory[  493] = 0;
        memory[  494] = 0;
        memory[  495] = 0;
        memory[  496] = 0;
        memory[  497] = 0;
        memory[  498] = 0;
        memory[  499] = 1;
        memory[  500] = 1;
        memory[  501] = 0;
        memory[  502] = 1;
        memory[  503] = 0;
        memory[  504] = 0;
        memory[  505] = 0;
        memory[  506] = 0;
        memory[  507] = 0;
        memory[  508] = 0;
        memory[  509] = 0;
        memory[  510] = 0;
        memory[  511] = 0;
        memory[  512] = 0;
        memory[  513] = 0;
        memory[  514] = 0;
        memory[  515] = 0;
        memory[  516] = 0;
        memory[  517] = 0;
        memory[  518] = 0;
        memory[  519] = 0;
        memory[  520] = 0;
        memory[  521] = 0;
        memory[  522] = 0;
        memory[  523] = 0;
        memory[  524] = 0;
        memory[  525] = 0;
        memory[  526] = 0;
        memory[  527] = 0;
        memory[  528] = 1;
        memory[  529] = 0;
        memory[  530] = 0;
        memory[  531] = 0;
        memory[  532] = 0;
        memory[  533] = 0;
        memory[  534] = 1;
        memory[  535] = 0;
        memory[  536] = 0;
        memory[  537] = 0;
        memory[  538] = 0;
        memory[  539] = 1;
        memory[  540] = 0;
        memory[  541] = 0;
        memory[  542] = 0;
        memory[  543] = 0;
        memory[  544] = 0;
        memory[  545] = 0;
        memory[  546] = 0;
        memory[  547] = 1;
        memory[  548] = 1;
        memory[  549] = 0;
        memory[  550] = 0;
        memory[  551] = 0;
        memory[  552] = 0;
        memory[  553] = 0;
        memory[  554] = 0;
        memory[  555] = 0;
        memory[  556] = 0;
        memory[  557] = 0;
        memory[  558] = 0;
        memory[  559] = 0;
        memory[  560] = 1;
        memory[  561] = 0;
        memory[  562] = 0;
        memory[  563] = 0;
        memory[  564] = 0;
        memory[  565] = 0;
        memory[  566] = 0;
        memory[  567] = 0;
        memory[  568] = 1;
        memory[  569] = 0;
        memory[  570] = 0;
        memory[  571] = 0;
        memory[  572] = 0;
        memory[  573] = 0;
        memory[  574] = 0;
        memory[  575] = 0;
        memory[  576] = 0;
        memory[  577] = 0;
        memory[  578] = 0;
        memory[  579] = 0;
        memory[  580] = 0;
        memory[  581] = 0;
        memory[  582] = 1;
        memory[  583] = 1;
        memory[  584] = 0;
        memory[  585] = 0;
        memory[  586] = 0;
        memory[  587] = 0;
        memory[  588] = 0;
        memory[  589] = 0;
        memory[  590] = 0;
        memory[  591] = 0;
        memory[  592] = 1;
        memory[  593] = 1;
        memory[  594] = 0;
        memory[  595] = 0;
        memory[  596] = 0;
        memory[  597] = 0;
        memory[  598] = 0;
        memory[  599] = 0;
        memory[  600] = 0;
        memory[  601] = 0;
        memory[  602] = 0;
        memory[  603] = 0;
        memory[  604] = 0;
        memory[  605] = 0;
        memory[  606] = 0;
        memory[  607] = 1;
        memory[  608] = 0;
        memory[  609] = 0;
        memory[  610] = 1;
        memory[  611] = 0;
        memory[  612] = 0;
        memory[  613] = 0;
        memory[  614] = 0;
        memory[  615] = 0;
        memory[  616] = 0;
        memory[  617] = 0;
        memory[  618] = 0;
        memory[  619] = 0;
        memory[  620] = 0;
        memory[  621] = 0;
        memory[  622] = 0;
        memory[  623] = 0;
        memory[  624] = 0;
        memory[  625] = 0;
        memory[  626] = 0;
        memory[  627] = 0;
        memory[  628] = 1;
        memory[  629] = 0;
        memory[  630] = 1;
        memory[  631] = 1;
        memory[  632] = 0;
        memory[  633] = 0;
        memory[  634] = 0;
        memory[  635] = 0;
        memory[  636] = 0;
        memory[  637] = 0;
        memory[  638] = 0;
        memory[  639] = 0;
        memory[  640] = 0;
        memory[  641] = 0;
        memory[  642] = 0;
        memory[  643] = 1;
        memory[  644] = 0;
        memory[  645] = 0;
        memory[  646] = 0;
        memory[  647] = 0;
        memory[  648] = 0;
        memory[  649] = 0;
        memory[  650] = 0;
        memory[  651] = 0;
        memory[  652] = 0;
        memory[  653] = 0;
        memory[  654] = 0;
        memory[  655] = 0;
        memory[  656] = 0;
        memory[  657] = 0;
        memory[  658] = 0;
        memory[  659] = 0;
        memory[  660] = 0;
        memory[  661] = 0;
        memory[  662] = 0;
        memory[  663] = 0;
        memory[  664] = 0;
        memory[  665] = 1;
        memory[  666] = 0;
        memory[  667] = 0;
        memory[  668] = 0;
        memory[  669] = 0;
        memory[  670] = 0;
        memory[  671] = 0;
        memory[  672] = 0;
        memory[  673] = 0;
        memory[  674] = 0;
        memory[  675] = 0;
        memory[  676] = 0;
        memory[  677] = 0;
        memory[  678] = 0;
        memory[  679] = 0;
        memory[  680] = 0;
        memory[  681] = 0;
        memory[  682] = 0;
        memory[  683] = 0;
        memory[  684] = 0;
        memory[  685] = 0;
        memory[  686] = 0;
        memory[  687] = 0;
        memory[  688] = 0;
        memory[  689] = 0;
        memory[  690] = 0;
        memory[  691] = 0;
        memory[  692] = 0;
        memory[  693] = 0;
        memory[  694] = 0;
        memory[  695] = 0;
        memory[  696] = 0;
        memory[  697] = 0;
        memory[  698] = 0;
        memory[  699] = 0;
        memory[  700] = 0;
        memory[  701] = 0;
        memory[  702] = 1;
        memory[  703] = 1;
        memory[  704] = 0;
        memory[  705] = 0;
        memory[  706] = 0;
        memory[  707] = 0;
        memory[  708] = 0;
        memory[  709] = 0;
        memory[  710] = 0;
        memory[  711] = 0;
        memory[  712] = 0;
        memory[  713] = 0;
        memory[  714] = 0;
        memory[  715] = 0;
        memory[  716] = 0;
        memory[  717] = 0;
        memory[  718] = 0;
        memory[  719] = 0;
        memory[  720] = 0;
        memory[  721] = 0;
        memory[  722] = 0;
        memory[  723] = 1;
        memory[  724] = 0;
        memory[  725] = 0;
        memory[  726] = 0;
        memory[  727] = 0;
        memory[  728] = 0;
        memory[  729] = 0;
        memory[  730] = 1;
        memory[  731] = 1;
        memory[  732] = 0;
        memory[  733] = 0;
        memory[  734] = 0;
        memory[  735] = 0;
        memory[  736] = 1;
        memory[  737] = 0;
        memory[  738] = 0;
        memory[  739] = 0;
        memory[  740] = 0;
        memory[  741] = 0;
        memory[  742] = 0;
        memory[  743] = 0;
        memory[  744] = 0;
        memory[  745] = 0;
        memory[  746] = 0;
        memory[  747] = 0;
        memory[  748] = 0;
        memory[  749] = 1;
        memory[  750] = 0;
        memory[  751] = 0;
        memory[  752] = 0;
        memory[  753] = 0;
        memory[  754] = 0;
        memory[  755] = 0;
        memory[  756] = 0;
        memory[  757] = 0;
        memory[  758] = 0;
        memory[  759] = 0;
        memory[  760] = 0;
        memory[  761] = 0;
        memory[  762] = 0;
        memory[  763] = 1;
        memory[  764] = 1;
        memory[  765] = 0;
        memory[  766] = 0;
        memory[  767] = 0;
        memory[  768] = 0;
        memory[  769] = 0;
        memory[  770] = 0;
        memory[  771] = 0;
        memory[  772] = 0;
        memory[  773] = 0;
        memory[  774] = 0;
        memory[  775] = 0;
        memory[  776] = 0;
        memory[  777] = 0;
        memory[  778] = 0;
        memory[  779] = 0;
        memory[  780] = 0;
        memory[  781] = 0;
        memory[  782] = 0;
        memory[  783] = 0;
        memory[  784] = 0;
        memory[  785] = 0;
        memory[  786] = 0;
        memory[  787] = 0;
        memory[  788] = 0;
        memory[  789] = 0;
        memory[  790] = 0;
        memory[  791] = 0;
        memory[  792] = 0;
        memory[  793] = 0;
        memory[  794] = 0;
        memory[  795] = 0;
        memory[  796] = 0;
        memory[  797] = 0;
        memory[  798] = 0;
        memory[  799] = 0;
        memory[  800] = 0;
        memory[  801] = 1;
        memory[  802] = 0;
        memory[  803] = 0;
        memory[  804] = 0;
        memory[  805] = 0;
        memory[  806] = 0;
        memory[  807] = 0;
        memory[  808] = 0;
        memory[  809] = 0;
        memory[  810] = 0;
        memory[  811] = 0;
        memory[  812] = 1;
        memory[  813] = 1;
        memory[  814] = 0;
        memory[  815] = 0;
        memory[  816] = 0;
        memory[  817] = 0;
        memory[  818] = 0;
        memory[  819] = 0;
        memory[  820] = 0;
        memory[  821] = 0;
        memory[  822] = 1;
        memory[  823] = 1;
        memory[  824] = 0;
        memory[  825] = 0;
        memory[  826] = 0;
        memory[  827] = 0;
        memory[  828] = 0;
        memory[  829] = 0;
        memory[  830] = 0;
        memory[  831] = 1;
        memory[  832] = 1;
        memory[  833] = 1;
        memory[  834] = 1;
        memory[  835] = 0;
        memory[  836] = 0;
        memory[  837] = 0;
        memory[  838] = 0;
        memory[  839] = 0;
        memory[  840] = 0;
        memory[  841] = 0;
        memory[  842] = 0;
        memory[  843] = 0;
        memory[  844] = 0;
        memory[  845] = 0;
        memory[  846] = 0;
        memory[  847] = 0;
        memory[  848] = 0;
        memory[  849] = 0;
        memory[  850] = 0;
        memory[  851] = 0;
        memory[  852] = 0;
        memory[  853] = 0;
        memory[  854] = 0;
        memory[  855] = 0;
        memory[  856] = 0;
        memory[  857] = 0;
        memory[  858] = 0;
        memory[  859] = 0;
        memory[  860] = 0;
        memory[  861] = 0;
        memory[  862] = 0;
        memory[  863] = 0;
        memory[  864] = 0;
        memory[  865] = 0;
        memory[  866] = 1;
        memory[  867] = 0;
        memory[  868] = 0;
        memory[  869] = 0;
        memory[  870] = 0;
        memory[  871] = 0;
        memory[  872] = 0;
        memory[  873] = 0;
        memory[  874] = 0;
        memory[  875] = 0;
        memory[  876] = 0;
        memory[  877] = 0;
        memory[  878] = 1;
        memory[  879] = 0;
        memory[  880] = 0;
        memory[  881] = 0;
        memory[  882] = 0;
        memory[  883] = 0;
        memory[  884] = 0;
        memory[  885] = 0;
        memory[  886] = 0;
        memory[  887] = 0;
        memory[  888] = 0;
        memory[  889] = 0;
        memory[  890] = 0;
        memory[  891] = 0;
        memory[  892] = 0;
        memory[  893] = 1;
        memory[  894] = 0;
        memory[  895] = 0;
        memory[  896] = 0;
        memory[  897] = 1;
        memory[  898] = 1;
        memory[  899] = 0;
        memory[  900] = 0;
        memory[  901] = 0;
        memory[  902] = 0;
        memory[  903] = 0;
        memory[  904] = 1;
        memory[  905] = 0;
        memory[  906] = 0;
        memory[  907] = 0;
        memory[  908] = 0;
        memory[  909] = 0;
        memory[  910] = 0;
        memory[  911] = 0;
        memory[  912] = 1;
        memory[  913] = 0;
        memory[  914] = 0;
        memory[  915] = 0;
        memory[  916] = 0;
        memory[  917] = 0;
        memory[  918] = 0;
        memory[  919] = 0;
        memory[  920] = 0;
        memory[  921] = 0;
        memory[  922] = 0;
        memory[  923] = 0;
        memory[  924] = 0;
        memory[  925] = 0;
        memory[  926] = 0;
        memory[  927] = 0;
        memory[  928] = 1;
        memory[  929] = 0;
        memory[  930] = 0;
        memory[  931] = 0;
        memory[  932] = 1;
        memory[  933] = 0;
        memory[  934] = 0;
        memory[  935] = 0;
        memory[  936] = 0;
        memory[  937] = 0;
        memory[  938] = 1;
        memory[  939] = 1;
        memory[  940] = 0;
        memory[  941] = 0;
        memory[  942] = 0;
        memory[  943] = 0;
        memory[  944] = 0;
        memory[  945] = 0;
        memory[  946] = 1;
        memory[  947] = 0;
        memory[  948] = 0;
        memory[  949] = 0;
        memory[  950] = 1;
        memory[  951] = 0;
        memory[  952] = 0;
        memory[  953] = 0;
        memory[  954] = 0;
        memory[  955] = 0;
        memory[  956] = 0;
        memory[  957] = 0;
        memory[  958] = 0;
        memory[  959] = 1;
        memory[  960] = 0;
        memory[  961] = 0;
        memory[  962] = 0;
        memory[  963] = 0;
        memory[  964] = 0;
        memory[  965] = 0;
        memory[  966] = 1;
        memory[  967] = 1;
        memory[  968] = 1;
        memory[  969] = 0;
        memory[  970] = 0;
        memory[  971] = 0;
        memory[  972] = 0;
        memory[  973] = 0;
        memory[  974] = 0;
        memory[  975] = 1;
        memory[  976] = 0;
        memory[  977] = 0;
        memory[  978] = 0;
        memory[  979] = 1;
        memory[  980] = 0;
        memory[  981] = 0;
        memory[  982] = 0;
        memory[  983] = 0;
        memory[  984] = 0;
        memory[  985] = 0;
        memory[  986] = 0;
        memory[  987] = 0;
        memory[  988] = 0;
        memory[  989] = 0;
        memory[  990] = 0;
        memory[  991] = 1;
        memory[  992] = 1;
        memory[  993] = 1;
        memory[  994] = 0;
        memory[  995] = 0;
        memory[  996] = 0;
        memory[  997] = 0;
        memory[  998] = 0;
        memory[  999] = 0;
        memory[ 1000] = 0;
        memory[ 1001] = 0;
        memory[ 1002] = 0;
        memory[ 1003] = 0;
        memory[ 1004] = 1;
        memory[ 1005] = 0;
        memory[ 1006] = 0;
        memory[ 1007] = 0;
        memory[ 1008] = 0;
        memory[ 1009] = 0;
        memory[ 1010] = 0;
        memory[ 1011] = 0;
        memory[ 1012] = 0;
        memory[ 1013] = 0;
        memory[ 1014] = 0;
        memory[ 1015] = 0;
        memory[ 1016] = 0;
        memory[ 1017] = 0;
        memory[ 1018] = 0;
        memory[ 1019] = 0;
        memory[ 1020] = 1;
        memory[ 1021] = 1;
        memory[ 1022] = 0;
        memory[ 1023] = 0;
        memory[ 1024] = 0;
        memory[ 1025] = 0;
        memory[ 1026] = 1;
        memory[ 1027] = 0;
        memory[ 1028] = 0;
        memory[ 1029] = 0;
        memory[ 1030] = 0;
        memory[ 1031] = 0;
        memory[ 1032] = 0;
        memory[ 1033] = 0;
        memory[ 1034] = 0;
        memory[ 1035] = 0;
        memory[ 1036] = 0;
        memory[ 1037] = 0;
        memory[ 1038] = 0;
        memory[ 1039] = 0;
        memory[ 1040] = 0;
        memory[ 1041] = 1;
        memory[ 1042] = 0;
        memory[ 1043] = 0;
        memory[ 1044] = 1;
        memory[ 1045] = 1;
        memory[ 1046] = 0;
        memory[ 1047] = 0;
        memory[ 1048] = 0;
        memory[ 1049] = 0;
        memory[ 1050] = 0;
        memory[ 1051] = 0;
        memory[ 1052] = 0;
        memory[ 1053] = 0;
        memory[ 1054] = 0;
        memory[ 1055] = 0;
        memory[ 1056] = 0;
        memory[ 1057] = 0;
        memory[ 1058] = 0;
        memory[ 1059] = 0;
        memory[ 1060] = 0;
        memory[ 1061] = 1;
        memory[ 1062] = 0;
        memory[ 1063] = 0;
        memory[ 1064] = 0;
        memory[ 1065] = 0;
        memory[ 1066] = 0;
        memory[ 1067] = 0;
        memory[ 1068] = 0;
        memory[ 1069] = 0;
        memory[ 1070] = 1;
        memory[ 1071] = 0;
        memory[ 1072] = 0;
        memory[ 1073] = 0;
        memory[ 1074] = 0;
        memory[ 1075] = 0;
        memory[ 1076] = 0;
        memory[ 1077] = 1;
        memory[ 1078] = 0;
        memory[ 1079] = 0;
        memory[ 1080] = 0;
        memory[ 1081] = 0;
        memory[ 1082] = 0;
        memory[ 1083] = 0;
        memory[ 1084] = 0;
        memory[ 1085] = 0;
        memory[ 1086] = 0;
        memory[ 1087] = 0;
        memory[ 1088] = 0;
        memory[ 1089] = 0;
        memory[ 1090] = 0;
        memory[ 1091] = 1;
        memory[ 1092] = 0;
        memory[ 1093] = 1;
        memory[ 1094] = 0;
        memory[ 1095] = 0;
        memory[ 1096] = 0;
        memory[ 1097] = 0;
        memory[ 1098] = 0;
        memory[ 1099] = 0;
        memory[ 1100] = 0;
        memory[ 1101] = 1;
        memory[ 1102] = 0;
        memory[ 1103] = 0;
        memory[ 1104] = 0;
        memory[ 1105] = 1;
        memory[ 1106] = 0;
        memory[ 1107] = 0;
        memory[ 1108] = 0;
        memory[ 1109] = 0;
        memory[ 1110] = 0;
        memory[ 1111] = 0;
        memory[ 1112] = 1;
        memory[ 1113] = 1;
        memory[ 1114] = 0;
        memory[ 1115] = 0;
        memory[ 1116] = 0;
        memory[ 1117] = 0;
        memory[ 1118] = 0;
        memory[ 1119] = 0;
        memory[ 1120] = 0;
        memory[ 1121] = 0;
        memory[ 1122] = 0;
        memory[ 1123] = 0;
        memory[ 1124] = 0;
        memory[ 1125] = 0;
        memory[ 1126] = 0;
        memory[ 1127] = 0;
        memory[ 1128] = 0;
        memory[ 1129] = 0;
        memory[ 1130] = 0;
        memory[ 1131] = 1;
        memory[ 1132] = 0;
        memory[ 1133] = 0;
        memory[ 1134] = 0;
        memory[ 1135] = 0;
        memory[ 1136] = 0;
        memory[ 1137] = 0;
        memory[ 1138] = 0;
        memory[ 1139] = 0;
        memory[ 1140] = 0;
        memory[ 1141] = 0;
        memory[ 1142] = 0;
        memory[ 1143] = 0;
        memory[ 1144] = 0;
        memory[ 1145] = 0;
        memory[ 1146] = 0;
        memory[ 1147] = 0;
        memory[ 1148] = 0;
        memory[ 1149] = 0;
        memory[ 1150] = 1;
        memory[ 1151] = 0;
        memory[ 1152] = 0;
        memory[ 1153] = 0;
        memory[ 1154] = 0;
        memory[ 1155] = 0;
        memory[ 1156] = 0;
        memory[ 1157] = 0;
        memory[ 1158] = 0;
        memory[ 1159] = 0;
        memory[ 1160] = 0;
        memory[ 1161] = 0;
        memory[ 1162] = 0;
        memory[ 1163] = 1;
        memory[ 1164] = 1;
        memory[ 1165] = 0;
        memory[ 1166] = 0;
        memory[ 1167] = 0;
        memory[ 1168] = 0;
        memory[ 1169] = 0;
        memory[ 1170] = 0;
        memory[ 1171] = 0;
        memory[ 1172] = 0;
        memory[ 1173] = 0;
        memory[ 1174] = 0;
        memory[ 1175] = 0;
        memory[ 1176] = 1;
        memory[ 1177] = 0;
        memory[ 1178] = 0;
        memory[ 1179] = 0;
        memory[ 1180] = 0;
        memory[ 1181] = 0;
        memory[ 1182] = 0;
        memory[ 1183] = 0;
        memory[ 1184] = 0;
        memory[ 1185] = 0;
        memory[ 1186] = 0;
        memory[ 1187] = 0;
        memory[ 1188] = 0;
        memory[ 1189] = 0;
        memory[ 1190] = 0;
        memory[ 1191] = 1;
        memory[ 1192] = 1;
        memory[ 1193] = 1;
        memory[ 1194] = 1;
        memory[ 1195] = 1;
        memory[ 1196] = 0;
        memory[ 1197] = 0;
        memory[ 1198] = 0;
        memory[ 1199] = 0;
        memory[ 1200] = 0;
        memory[ 1201] = 0;
        memory[ 1202] = 0;
        memory[ 1203] = 0;
        memory[ 1204] = 1;
        memory[ 1205] = 0;
        memory[ 1206] = 0;
        memory[ 1207] = 0;
        memory[ 1208] = 1;
        memory[ 1209] = 1;
        memory[ 1210] = 0;
        memory[ 1211] = 0;
        memory[ 1212] = 0;
        memory[ 1213] = 0;
        memory[ 1214] = 0;
        memory[ 1215] = 0;
        memory[ 1216] = 0;
        memory[ 1217] = 0;
        memory[ 1218] = 1;
        memory[ 1219] = 0;
        memory[ 1220] = 0;
        memory[ 1221] = 1;
        memory[ 1222] = 1;
        memory[ 1223] = 0;
        memory[ 1224] = 0;
        memory[ 1225] = 0;
        memory[ 1226] = 0;
        memory[ 1227] = 0;
        memory[ 1228] = 0;
        memory[ 1229] = 0;
        memory[ 1230] = 0;
        memory[ 1231] = 0;
        memory[ 1232] = 0;
        memory[ 1233] = 0;
        memory[ 1234] = 0;
        memory[ 1235] = 0;
        memory[ 1236] = 0;
        memory[ 1237] = 1;
        memory[ 1238] = 0;
        memory[ 1239] = 0;
        memory[ 1240] = 0;
        memory[ 1241] = 0;
        memory[ 1242] = 0;
        memory[ 1243] = 0;
        memory[ 1244] = 0;
        memory[ 1245] = 0;
        memory[ 1246] = 0;
        memory[ 1247] = 0;
        memory[ 1248] = 0;
        memory[ 1249] = 0;
        memory[ 1250] = 0;
        memory[ 1251] = 0;
        memory[ 1252] = 0;
        memory[ 1253] = 0;
        memory[ 1254] = 0;
        memory[ 1255] = 1;
        memory[ 1256] = 0;
        memory[ 1257] = 0;
        memory[ 1258] = 0;
        memory[ 1259] = 0;
        memory[ 1260] = 0;
        memory[ 1261] = 0;
        memory[ 1262] = 0;
        memory[ 1263] = 0;
        memory[ 1264] = 0;
        memory[ 1265] = 0;
        memory[ 1266] = 0;
        memory[ 1267] = 0;
        memory[ 1268] = 0;
        memory[ 1269] = 0;
        memory[ 1270] = 0;
        memory[ 1271] = 0;
        memory[ 1272] = 0;
        memory[ 1273] = 0;
        memory[ 1274] = 0;
        memory[ 1275] = 0;
        memory[ 1276] = 0;
        memory[ 1277] = 0;
        memory[ 1278] = 0;
        memory[ 1279] = 0;
        memory[ 1280] = 0;
        memory[ 1281] = 1;
        memory[ 1282] = 1;
        memory[ 1283] = 0;
        memory[ 1284] = 0;
        memory[ 1285] = 0;
        memory[ 1286] = 0;
        memory[ 1287] = 0;
        memory[ 1288] = 0;
        memory[ 1289] = 0;
        memory[ 1290] = 0;
        memory[ 1291] = 0;
        memory[ 1292] = 0;
        memory[ 1293] = 1;
        memory[ 1294] = 1;
        memory[ 1295] = 0;
        memory[ 1296] = 0;
        memory[ 1297] = 0;
        memory[ 1298] = 0;
        memory[ 1299] = 0;
        memory[ 1300] = 0;
        memory[ 1301] = 0;
        memory[ 1302] = 0;
        memory[ 1303] = 0;
        memory[ 1304] = 0;
        memory[ 1305] = 0;
        memory[ 1306] = 0;
        memory[ 1307] = 0;
        memory[ 1308] = 0;
        memory[ 1309] = 0;
        memory[ 1310] = 1;
        memory[ 1311] = 0;
        memory[ 1312] = 0;
        memory[ 1313] = 0;
        memory[ 1314] = 0;
        memory[ 1315] = 0;
        memory[ 1316] = 0;
        memory[ 1317] = 0;
        memory[ 1318] = 0;
        memory[ 1319] = 0;
        memory[ 1320] = 0;
        memory[ 1321] = 0;
        memory[ 1322] = 0;
        memory[ 1323] = 0;
        memory[ 1324] = 0;
        memory[ 1325] = 0;
        memory[ 1326] = 0;
        memory[ 1327] = 1;
        memory[ 1328] = 0;
        memory[ 1329] = 0;
        memory[ 1330] = 1;
        memory[ 1331] = 0;
        memory[ 1332] = 0;
        memory[ 1333] = 0;
        memory[ 1334] = 0;
        memory[ 1335] = 0;
        memory[ 1336] = 0;
        memory[ 1337] = 0;
        memory[ 1338] = 0;
        memory[ 1339] = 0;
        memory[ 1340] = 0;
        memory[ 1341] = 0;
        memory[ 1342] = 0;
        memory[ 1343] = 1;
        memory[ 1344] = 0;
        memory[ 1345] = 0;
        memory[ 1346] = 0;
        memory[ 1347] = 0;
        memory[ 1348] = 0;
        memory[ 1349] = 0;
        memory[ 1350] = 0;
        memory[ 1351] = 0;
        memory[ 1352] = 0;
        memory[ 1353] = 0;
        memory[ 1354] = 0;
        memory[ 1355] = 0;
        memory[ 1356] = 0;
        memory[ 1357] = 0;
        memory[ 1358] = 0;
        memory[ 1359] = 0;
        memory[ 1360] = 0;
        memory[ 1361] = 0;
        memory[ 1362] = 0;
        memory[ 1363] = 0;
        memory[ 1364] = 0;
        memory[ 1365] = 0;
        memory[ 1366] = 0;
        memory[ 1367] = 0;
        memory[ 1368] = 0;
        memory[ 1369] = 0;
        memory[ 1370] = 0;
        memory[ 1371] = 1;
        memory[ 1372] = 0;
        memory[ 1373] = 1;
        memory[ 1374] = 0;
        memory[ 1375] = 0;
        memory[ 1376] = 0;
        memory[ 1377] = 0;
        memory[ 1378] = 0;
        memory[ 1379] = 0;
        memory[ 1380] = 0;
        memory[ 1381] = 0;
        memory[ 1382] = 0;
        memory[ 1383] = 0;
        memory[ 1384] = 0;
        memory[ 1385] = 0;
        memory[ 1386] = 0;
        memory[ 1387] = 1;
        memory[ 1388] = 1;
        memory[ 1389] = 0;
        memory[ 1390] = 0;
        memory[ 1391] = 0;
        memory[ 1392] = 0;
        memory[ 1393] = 0;
        memory[ 1394] = 1;
        memory[ 1395] = 1;
        memory[ 1396] = 0;
        memory[ 1397] = 0;
        memory[ 1398] = 0;
        memory[ 1399] = 0;
        memory[ 1400] = 0;
        memory[ 1401] = 0;
        memory[ 1402] = 0;
        memory[ 1403] = 0;
        memory[ 1404] = 0;
        memory[ 1405] = 1;
        memory[ 1406] = 1;
        memory[ 1407] = 0;
        memory[ 1408] = 0;
        memory[ 1409] = 0;
        memory[ 1410] = 0;
        memory[ 1411] = 0;
        memory[ 1412] = 0;
        memory[ 1413] = 0;
        memory[ 1414] = 0;
        memory[ 1415] = 0;
        memory[ 1416] = 0;
        memory[ 1417] = 0;
        memory[ 1418] = 0;
        memory[ 1419] = 0;
        memory[ 1420] = 0;
        memory[ 1421] = 0;
        memory[ 1422] = 0;
        memory[ 1423] = 0;
        memory[ 1424] = 0;
        memory[ 1425] = 0;
        memory[ 1426] = 0;
        memory[ 1427] = 1;
        memory[ 1428] = 0;
        memory[ 1429] = 0;
        memory[ 1430] = 0;
        memory[ 1431] = 0;
        memory[ 1432] = 0;
        memory[ 1433] = 0;
        memory[ 1434] = 0;
        memory[ 1435] = 1;
        memory[ 1436] = 0;
        memory[ 1437] = 0;
        memory[ 1438] = 0;
        memory[ 1439] = 0;
        memory[ 1440] = 0;
        memory[ 1441] = 0;
        memory[ 1442] = 0;
        memory[ 1443] = 0;
        memory[ 1444] = 0;
        memory[ 1445] = 0;
        memory[ 1446] = 0;
        memory[ 1447] = 0;
        memory[ 1448] = 0;
        memory[ 1449] = 0;
        memory[ 1450] = 0;
        memory[ 1451] = 0;
        memory[ 1452] = 0;
        memory[ 1453] = 0;
        memory[ 1454] = 0;
        memory[ 1455] = 1;
        memory[ 1456] = 0;
        memory[ 1457] = 0;
        memory[ 1458] = 0;
        memory[ 1459] = 0;
        memory[ 1460] = 1;
        memory[ 1461] = 0;
        memory[ 1462] = 0;
        memory[ 1463] = 0;
        memory[ 1464] = 0;
        memory[ 1465] = 0;
        memory[ 1466] = 0;
        memory[ 1467] = 0;
        memory[ 1468] = 0;
        memory[ 1469] = 0;
        memory[ 1470] = 0;
        memory[ 1471] = 1;
        memory[ 1472] = 0;
        memory[ 1473] = 0;
        memory[ 1474] = 0;
        memory[ 1475] = 0;
        memory[ 1476] = 0;
        memory[ 1477] = 0;
        memory[ 1478] = 0;
        memory[ 1479] = 0;
        memory[ 1480] = 0;
        memory[ 1481] = 0;
        memory[ 1482] = 0;
        memory[ 1483] = 0;
        memory[ 1484] = 0;
        memory[ 1485] = 0;
        memory[ 1486] = 0;
        memory[ 1487] = 0;
        memory[ 1488] = 0;
        memory[ 1489] = 0;
        memory[ 1490] = 0;
        memory[ 1491] = 0;
        memory[ 1492] = 0;
        memory[ 1493] = 0;
        memory[ 1494] = 0;
        memory[ 1495] = 0;
        memory[ 1496] = 0;
        memory[ 1497] = 1;
        memory[ 1498] = 0;
        memory[ 1499] = 0;
        memory[ 1500] = 0;
        memory[ 1501] = 0;
        memory[ 1502] = 0;
        memory[ 1503] = 0;
        memory[ 1504] = 0;
        memory[ 1505] = 0;
        memory[ 1506] = 0;
        memory[ 1507] = 0;
        memory[ 1508] = 0;
        memory[ 1509] = 0;
        memory[ 1510] = 0;
        memory[ 1511] = 1;
        memory[ 1512] = 0;
        memory[ 1513] = 0;
        memory[ 1514] = 0;
        memory[ 1515] = 0;
        memory[ 1516] = 0;
        memory[ 1517] = 0;
        memory[ 1518] = 1;
        memory[ 1519] = 1;
        memory[ 1520] = 0;
        memory[ 1521] = 0;
        memory[ 1522] = 0;
        memory[ 1523] = 0;
        memory[ 1524] = 0;
        memory[ 1525] = 1;
        memory[ 1526] = 1;
        memory[ 1527] = 0;
        memory[ 1528] = 0;
        memory[ 1529] = 0;
        memory[ 1530] = 0;
        memory[ 1531] = 0;
        memory[ 1532] = 0;
        memory[ 1533] = 0;
        memory[ 1534] = 0;
        memory[ 1535] = 0;
        memory[ 1536] = 0;
        memory[ 1537] = 0;
        memory[ 1538] = 0;
        memory[ 1539] = 0;
        memory[ 1540] = 0;
        memory[ 1541] = 0;
        memory[ 1542] = 0;
        memory[ 1543] = 0;
        memory[ 1544] = 0;
        memory[ 1545] = 0;
        memory[ 1546] = 0;
        memory[ 1547] = 0;
        memory[ 1548] = 0;
        memory[ 1549] = 0;
        memory[ 1550] = 1;
        memory[ 1551] = 0;
        memory[ 1552] = 0;
        memory[ 1553] = 0;
        memory[ 1554] = 1;
        memory[ 1555] = 1;
        memory[ 1556] = 0;
        memory[ 1557] = 0;
        memory[ 1558] = 0;
        memory[ 1559] = 0;
        memory[ 1560] = 0;
        memory[ 1561] = 0;
        memory[ 1562] = 0;
        memory[ 1563] = 0;
        memory[ 1564] = 0;
        memory[ 1565] = 0;
        memory[ 1566] = 0;
        memory[ 1567] = 1;
        memory[ 1568] = 0;
        memory[ 1569] = 0;
        memory[ 1570] = 0;
        memory[ 1571] = 0;
        memory[ 1572] = 0;
        memory[ 1573] = 0;
        memory[ 1574] = 0;
        memory[ 1575] = 1;
        memory[ 1576] = 1;
        memory[ 1577] = 0;
        memory[ 1578] = 0;
        memory[ 1579] = 0;
        memory[ 1580] = 0;
        memory[ 1581] = 0;
        memory[ 1582] = 0;
        memory[ 1583] = 0;
        memory[ 1584] = 0;
        memory[ 1585] = 0;
        memory[ 1586] = 0;
        memory[ 1587] = 0;
        memory[ 1588] = 0;
        memory[ 1589] = 0;
        memory[ 1590] = 0;
        memory[ 1591] = 0;
        memory[ 1592] = 0;
        memory[ 1593] = 0;
        memory[ 1594] = 0;
        memory[ 1595] = 0;
        memory[ 1596] = 0;
        memory[ 1597] = 0;
        memory[ 1598] = 0;
        memory[ 1599] = 0;
        memory[ 1600] = 0;
        memory[ 1601] = 0;
        memory[ 1602] = 0;
        memory[ 1603] = 0;
        memory[ 1604] = 0;
        memory[ 1605] = 1;
        memory[ 1606] = 1;
        memory[ 1607] = 0;
        memory[ 1608] = 0;
        memory[ 1609] = 0;
        memory[ 1610] = 1;
        memory[ 1611] = 0;
        memory[ 1612] = 0;
        memory[ 1613] = 0;
        memory[ 1614] = 0;
        memory[ 1615] = 0;
        memory[ 1616] = 1;
        memory[ 1617] = 0;
        memory[ 1618] = 0;
        memory[ 1619] = 0;
        memory[ 1620] = 0;
        memory[ 1621] = 0;
        memory[ 1622] = 0;
        memory[ 1623] = 0;
        memory[ 1624] = 0;
        memory[ 1625] = 0;
        memory[ 1626] = 0;
        memory[ 1627] = 0;
        memory[ 1628] = 0;
        memory[ 1629] = 0;
        memory[ 1630] = 0;
        memory[ 1631] = 0;
        memory[ 1632] = 0;
        memory[ 1633] = 0;
        memory[ 1634] = 0;
        memory[ 1635] = 0;
        memory[ 1636] = 0;
        memory[ 1637] = 0;
        memory[ 1638] = 0;
        memory[ 1639] = 1;
        memory[ 1640] = 0;
        memory[ 1641] = 0;
        memory[ 1642] = 0;
        memory[ 1643] = 0;
        memory[ 1644] = 0;
        memory[ 1645] = 0;
        memory[ 1646] = 0;
        memory[ 1647] = 1;
        memory[ 1648] = 0;
        memory[ 1649] = 0;
        memory[ 1650] = 0;
        memory[ 1651] = 0;
        memory[ 1652] = 0;
        memory[ 1653] = 0;
        memory[ 1654] = 1;
        memory[ 1655] = 1;
        memory[ 1656] = 0;
        memory[ 1657] = 0;
        memory[ 1658] = 0;
        memory[ 1659] = 0;
        memory[ 1660] = 0;
        memory[ 1661] = 0;
        memory[ 1662] = 0;
        memory[ 1663] = 0;
        memory[ 1664] = 0;
        memory[ 1665] = 0;
        memory[ 1666] = 0;
        memory[ 1667] = 0;
        memory[ 1668] = 0;
        memory[ 1669] = 0;
        memory[ 1670] = 0;
        memory[ 1671] = 0;
        memory[ 1672] = 0;
        memory[ 1673] = 0;
        memory[ 1674] = 0;
        memory[ 1675] = 0;
        memory[ 1676] = 0;
        memory[ 1677] = 0;
        memory[ 1678] = 0;
        memory[ 1679] = 0;
        memory[ 1680] = 0;
        memory[ 1681] = 0;
        memory[ 1682] = 0;
        memory[ 1683] = 0;
        memory[ 1684] = 0;
        memory[ 1685] = 0;
        memory[ 1686] = 0;
        memory[ 1687] = 1;
        memory[ 1688] = 0;
        memory[ 1689] = 1;
        memory[ 1690] = 0;
        memory[ 1691] = 0;
        memory[ 1692] = 0;
        memory[ 1693] = 0;
        memory[ 1694] = 1;
        memory[ 1695] = 0;
        memory[ 1696] = 0;
        memory[ 1697] = 0;
        memory[ 1698] = 0;
        memory[ 1699] = 0;
        memory[ 1700] = 0;
        memory[ 1701] = 0;
        memory[ 1702] = 0;
        memory[ 1703] = 0;
        memory[ 1704] = 0;
        memory[ 1705] = 1;
        memory[ 1706] = 1;
        memory[ 1707] = 0;
        memory[ 1708] = 0;
        memory[ 1709] = 0;
        memory[ 1710] = 0;
        memory[ 1711] = 1;
        memory[ 1712] = 1;
        memory[ 1713] = 0;
        memory[ 1714] = 1;
        memory[ 1715] = 0;
        memory[ 1716] = 0;
        memory[ 1717] = 0;
        memory[ 1718] = 0;
        memory[ 1719] = 0;
        memory[ 1720] = 0;
        memory[ 1721] = 0;
        memory[ 1722] = 0;
        memory[ 1723] = 0;
        memory[ 1724] = 0;
        memory[ 1725] = 0;
        memory[ 1726] = 0;
        memory[ 1727] = 0;
        memory[ 1728] = 0;
        memory[ 1729] = 0;
        memory[ 1730] = 0;
        memory[ 1731] = 0;
        memory[ 1732] = 1;
        memory[ 1733] = 0;
        memory[ 1734] = 0;
        memory[ 1735] = 0;
        memory[ 1736] = 0;
        memory[ 1737] = 0;
        memory[ 1738] = 0;
        memory[ 1739] = 1;
        memory[ 1740] = 0;
        memory[ 1741] = 0;
        memory[ 1742] = 0;
        memory[ 1743] = 0;
        memory[ 1744] = 1;
        memory[ 1745] = 0;
        memory[ 1746] = 0;
        memory[ 1747] = 0;
        memory[ 1748] = 0;
        memory[ 1749] = 0;
        memory[ 1750] = 0;
        memory[ 1751] = 0;
        memory[ 1752] = 0;
        memory[ 1753] = 0;
        memory[ 1754] = 0;
        memory[ 1755] = 0;
        memory[ 1756] = 0;
        memory[ 1757] = 1;
        memory[ 1758] = 0;
        memory[ 1759] = 0;
        memory[ 1760] = 0;
        memory[ 1761] = 0;
        memory[ 1762] = 0;
        memory[ 1763] = 0;
        memory[ 1764] = 0;
        memory[ 1765] = 0;
        memory[ 1766] = 0;
        memory[ 1767] = 0;
        memory[ 1768] = 0;
        memory[ 1769] = 0;
        memory[ 1770] = 0;
        memory[ 1771] = 0;
        memory[ 1772] = 0;
        memory[ 1773] = 0;
        memory[ 1774] = 0;
        memory[ 1775] = 1;
        memory[ 1776] = 0;
        memory[ 1777] = 0;
        memory[ 1778] = 0;
        memory[ 1779] = 1;
        memory[ 1780] = 1;
        memory[ 1781] = 0;
        memory[ 1782] = 0;
        memory[ 1783] = 0;
        memory[ 1784] = 0;
        memory[ 1785] = 0;
        memory[ 1786] = 0;
        memory[ 1787] = 0;
        memory[ 1788] = 1;
        memory[ 1789] = 1;
        memory[ 1790] = 1;
        memory[ 1791] = 0;
        memory[ 1792] = 0;
        memory[ 1793] = 1;
        memory[ 1794] = 0;
        memory[ 1795] = 1;
        memory[ 1796] = 1;
        memory[ 1797] = 0;
        memory[ 1798] = 0;
        memory[ 1799] = 0;
        memory[ 1800] = 0;
        memory[ 1801] = 0;
        memory[ 1802] = 1;
        memory[ 1803] = 0;
        memory[ 1804] = 0;
        memory[ 1805] = 0;
        memory[ 1806] = 0;
        memory[ 1807] = 0;
        memory[ 1808] = 0;
        memory[ 1809] = 0;
        memory[ 1810] = 0;
        memory[ 1811] = 0;
        memory[ 1812] = 0;
        memory[ 1813] = 0;
        memory[ 1814] = 0;
        memory[ 1815] = 0;
        memory[ 1816] = 0;
        memory[ 1817] = 0;
        memory[ 1818] = 1;
        memory[ 1819] = 0;
        memory[ 1820] = 0;
        memory[ 1821] = 0;
        memory[ 1822] = 0;
        memory[ 1823] = 0;
        memory[ 1824] = 0;
        memory[ 1825] = 0;
        memory[ 1826] = 0;
        memory[ 1827] = 0;
        memory[ 1828] = 0;
        memory[ 1829] = 0;
        memory[ 1830] = 0;
        memory[ 1831] = 0;
        memory[ 1832] = 0;
        memory[ 1833] = 0;
        memory[ 1834] = 0;
        memory[ 1835] = 0;
        memory[ 1836] = 0;
        memory[ 1837] = 0;
        memory[ 1838] = 0;
        memory[ 1839] = 1;
        memory[ 1840] = 0;
        memory[ 1841] = 0;
        memory[ 1842] = 0;
        memory[ 1843] = 0;
        memory[ 1844] = 0;
        memory[ 1845] = 0;
        memory[ 1846] = 0;
        memory[ 1847] = 0;
        memory[ 1848] = 1;
        memory[ 1849] = 0;
        memory[ 1850] = 0;
        memory[ 1851] = 0;
        memory[ 1852] = 0;
        memory[ 1853] = 0;
        memory[ 1854] = 0;
        memory[ 1855] = 0;
        memory[ 1856] = 0;
        memory[ 1857] = 0;
        memory[ 1858] = 0;
        memory[ 1859] = 0;
        memory[ 1860] = 0;
        memory[ 1861] = 0;
        memory[ 1862] = 0;
        memory[ 1863] = 0;
        memory[ 1864] = 0;
        memory[ 1865] = 0;
        memory[ 1866] = 0;
        memory[ 1867] = 0;
        memory[ 1868] = 0;
        memory[ 1869] = 0;
        memory[ 1870] = 0;
        memory[ 1871] = 0;
        memory[ 1872] = 1;
        memory[ 1873] = 1;
        memory[ 1874] = 0;
        memory[ 1875] = 1;
        memory[ 1876] = 1;
        memory[ 1877] = 1;
        memory[ 1878] = 0;
        memory[ 1879] = 1;
        memory[ 1880] = 0;
        memory[ 1881] = 0;
        memory[ 1882] = 0;
        memory[ 1883] = 0;
        memory[ 1884] = 0;
        memory[ 1885] = 0;
        memory[ 1886] = 0;
        memory[ 1887] = 0;
        memory[ 1888] = 0;
        memory[ 1889] = 0;
        memory[ 1890] = 1;
        memory[ 1891] = 1;
        memory[ 1892] = 0;
        memory[ 1893] = 0;
        memory[ 1894] = 0;
        memory[ 1895] = 0;
        memory[ 1896] = 0;
        memory[ 1897] = 0;
        memory[ 1898] = 0;
        memory[ 1899] = 0;
        memory[ 1900] = 0;
        memory[ 1901] = 0;
        memory[ 1902] = 0;
        memory[ 1903] = 0;
        memory[ 1904] = 0;
        memory[ 1905] = 0;
        memory[ 1906] = 0;
        memory[ 1907] = 0;
        memory[ 1908] = 0;
        memory[ 1909] = 0;
        memory[ 1910] = 0;
        memory[ 1911] = 0;
        memory[ 1912] = 0;
        memory[ 1913] = 0;
        memory[ 1914] = 0;
        memory[ 1915] = 0;
        memory[ 1916] = 0;
        memory[ 1917] = 0;
        memory[ 1918] = 0;
        memory[ 1919] = 0;
        memory[ 1920] = 0;
        memory[ 1921] = 0;
        memory[ 1922] = 0;
        memory[ 1923] = 0;
        memory[ 1924] = 0;
        memory[ 1925] = 0;
        memory[ 1926] = 0;
        memory[ 1927] = 0;
        memory[ 1928] = 0;
        memory[ 1929] = 0;
        memory[ 1930] = 0;
        memory[ 1931] = 0;
        memory[ 1932] = 0;
        memory[ 1933] = 0;
        memory[ 1934] = 0;
        memory[ 1935] = 0;
        memory[ 1936] = 0;
        memory[ 1937] = 0;
        memory[ 1938] = 0;
        memory[ 1939] = 0;
        memory[ 1940] = 0;
        memory[ 1941] = 0;
        memory[ 1942] = 0;
        memory[ 1943] = 0;
        memory[ 1944] = 0;
        memory[ 1945] = 0;
        memory[ 1946] = 1;
        memory[ 1947] = 0;
        memory[ 1948] = 0;
        memory[ 1949] = 0;
        memory[ 1950] = 0;
        memory[ 1951] = 0;
        memory[ 1952] = 0;
        memory[ 1953] = 0;
        memory[ 1954] = 0;
        memory[ 1955] = 0;
        memory[ 1956] = 0;
        memory[ 1957] = 0;
        memory[ 1958] = 0;
        memory[ 1959] = 1;
        memory[ 1960] = 0;
        memory[ 1961] = 0;
        memory[ 1962] = 1;
        memory[ 1963] = 0;
        memory[ 1964] = 0;
        memory[ 1965] = 1;
        memory[ 1966] = 0;
        memory[ 1967] = 0;
        memory[ 1968] = 0;
        memory[ 1969] = 1;
        memory[ 1970] = 0;
        memory[ 1971] = 0;
        memory[ 1972] = 0;
        memory[ 1973] = 0;
        memory[ 1974] = 0;
        memory[ 1975] = 0;
        memory[ 1976] = 0;
        memory[ 1977] = 0;
        memory[ 1978] = 0;
        memory[ 1979] = 0;
        memory[ 1980] = 0;
        memory[ 1981] = 0;
        memory[ 1982] = 0;
        memory[ 1983] = 0;
        memory[ 1984] = 0;
        memory[ 1985] = 0;
        memory[ 1986] = 0;
        memory[ 1987] = 0;
        memory[ 1988] = 0;
        memory[ 1989] = 0;
        memory[ 1990] = 0;
        memory[ 1991] = 0;
        memory[ 1992] = 0;
        memory[ 1993] = 0;
        memory[ 1994] = 0;
        memory[ 1995] = 0;
        memory[ 1996] = 0;
        memory[ 1997] = 0;
        memory[ 1998] = 0;
        memory[ 1999] = 0;
        memory[ 2000] = 0;
        memory[ 2001] = 0;
        memory[ 2002] = 0;
        memory[ 2003] = 0;
        memory[ 2004] = 0;
        memory[ 2005] = 0;
        memory[ 2006] = 0;
        memory[ 2007] = 0;
        memory[ 2008] = 0;
        memory[ 2009] = 0;
        memory[ 2010] = 0;
        memory[ 2011] = 0;
        memory[ 2012] = 0;
        memory[ 2013] = 0;
        memory[ 2014] = 0;
        memory[ 2015] = 0;
        memory[ 2016] = 0;
        memory[ 2017] = 0;
        memory[ 2018] = 0;
        memory[ 2019] = 0;
        memory[ 2020] = 0;
        memory[ 2021] = 0;
        memory[ 2022] = 0;
        memory[ 2023] = 0;
        memory[ 2024] = 0;
        memory[ 2025] = 0;
        memory[ 2026] = 0;
        memory[ 2027] = 0;
        memory[ 2028] = 0;
        memory[ 2029] = 0;
        memory[ 2030] = 0;
        memory[ 2031] = 0;
        memory[ 2032] = 0;
        memory[ 2033] = 0;
        memory[ 2034] = 0;
        memory[ 2035] = 0;
        memory[ 2036] = 0;
        memory[ 2037] = 0;
        memory[ 2038] = 0;
        memory[ 2039] = 0;
        memory[ 2040] = 0;
        memory[ 2041] = 0;
        memory[ 2042] = 0;
        memory[ 2043] = 0;
        memory[ 2044] = 0;
        memory[ 2045] = 0;
        memory[ 2046] = 0;
        memory[ 2047] = 0;
        memory[ 2048] = 1;
        memory[ 2049] = 0;
        memory[ 2050] = 0;
        memory[ 2051] = 0;
        memory[ 2052] = 0;
        memory[ 2053] = 0;
        memory[ 2054] = 0;
        memory[ 2055] = 0;
        memory[ 2056] = 0;
        memory[ 2057] = 0;
        memory[ 2058] = 0;
        memory[ 2059] = 0;
        memory[ 2060] = 1;
        memory[ 2061] = 0;
        memory[ 2062] = 0;
        memory[ 2063] = 0;
        memory[ 2064] = 0;
        memory[ 2065] = 0;
        memory[ 2066] = 0;
        memory[ 2067] = 0;
        memory[ 2068] = 0;
        memory[ 2069] = 0;
        memory[ 2070] = 0;
        memory[ 2071] = 0;
        memory[ 2072] = 0;
        memory[ 2073] = 0;
        memory[ 2074] = 0;
        memory[ 2075] = 0;
        memory[ 2076] = 0;
        memory[ 2077] = 0;
        memory[ 2078] = 0;
        memory[ 2079] = 0;
        memory[ 2080] = 0;
        memory[ 2081] = 0;
        memory[ 2082] = 0;
        memory[ 2083] = 0;
        memory[ 2084] = 0;
        memory[ 2085] = 0;
        memory[ 2086] = 1;
        memory[ 2087] = 0;
        memory[ 2088] = 0;
        memory[ 2089] = 0;
        memory[ 2090] = 0;
        memory[ 2091] = 0;
        memory[ 2092] = 1;
        memory[ 2093] = 0;
        memory[ 2094] = 0;
        memory[ 2095] = 0;
        memory[ 2096] = 0;
        memory[ 2097] = 0;
        memory[ 2098] = 0;
        memory[ 2099] = 0;
        memory[ 2100] = 0;
        memory[ 2101] = 0;
        memory[ 2102] = 0;
        memory[ 2103] = 0;
        memory[ 2104] = 0;
        memory[ 2105] = 0;
        memory[ 2106] = 0;
        memory[ 2107] = 0;
        memory[ 2108] = 0;
        memory[ 2109] = 0;
        memory[ 2110] = 0;
        memory[ 2111] = 0;
        memory[ 2112] = 0;
        memory[ 2113] = 0;
        memory[ 2114] = 0;
        memory[ 2115] = 0;
        memory[ 2116] = 0;
        memory[ 2117] = 0;
        memory[ 2118] = 0;
        memory[ 2119] = 0;
        memory[ 2120] = 0;
        memory[ 2121] = 0;
        memory[ 2122] = 0;
        memory[ 2123] = 0;
        memory[ 2124] = 0;
        memory[ 2125] = 0;
        memory[ 2126] = 0;
        memory[ 2127] = 0;
        memory[ 2128] = 0;
        memory[ 2129] = 0;
        memory[ 2130] = 0;
        memory[ 2131] = 0;
        memory[ 2132] = 0;
        memory[ 2133] = 0;
        memory[ 2134] = 0;
        memory[ 2135] = 0;
        memory[ 2136] = 0;
        memory[ 2137] = 0;
        memory[ 2138] = 0;
        memory[ 2139] = 0;
        memory[ 2140] = 0;
        memory[ 2141] = 1;
        memory[ 2142] = 1;
        memory[ 2143] = 0;
        memory[ 2144] = 0;
        memory[ 2145] = 0;
        memory[ 2146] = 0;
        memory[ 2147] = 0;
        memory[ 2148] = 0;
        memory[ 2149] = 1;
        memory[ 2150] = 1;
        memory[ 2151] = 0;
        memory[ 2152] = 0;
        memory[ 2153] = 0;
        memory[ 2154] = 0;
        memory[ 2155] = 0;
        memory[ 2156] = 0;
        memory[ 2157] = 0;
        memory[ 2158] = 1;
        memory[ 2159] = 0;
        memory[ 2160] = 0;
        memory[ 2161] = 0;
        memory[ 2162] = 0;
        memory[ 2163] = 0;
        memory[ 2164] = 0;
        memory[ 2165] = 0;
        memory[ 2166] = 0;
        memory[ 2167] = 0;
        memory[ 2168] = 0;
        memory[ 2169] = 0;
        memory[ 2170] = 0;
        memory[ 2171] = 1;
        memory[ 2172] = 1;
        memory[ 2173] = 0;
        memory[ 2174] = 0;
        memory[ 2175] = 0;
        memory[ 2176] = 0;
        memory[ 2177] = 0;
        memory[ 2178] = 0;
        memory[ 2179] = 0;
        memory[ 2180] = 0;
        memory[ 2181] = 0;
        memory[ 2182] = 0;
        memory[ 2183] = 0;
        memory[ 2184] = 0;
        memory[ 2185] = 0;
        memory[ 2186] = 0;
        memory[ 2187] = 0;
        memory[ 2188] = 0;
        memory[ 2189] = 0;
        memory[ 2190] = 0;
        memory[ 2191] = 0;
        memory[ 2192] = 0;
        memory[ 2193] = 0;
        memory[ 2194] = 0;
        memory[ 2195] = 0;
        memory[ 2196] = 0;
        memory[ 2197] = 0;
        memory[ 2198] = 0;
        memory[ 2199] = 0;
        memory[ 2200] = 0;
        memory[ 2201] = 0;
        memory[ 2202] = 0;
        memory[ 2203] = 0;
        memory[ 2204] = 0;
        memory[ 2205] = 0;
        memory[ 2206] = 0;
        memory[ 2207] = 0;
        memory[ 2208] = 0;
        memory[ 2209] = 0;
        memory[ 2210] = 0;
        memory[ 2211] = 0;
        memory[ 2212] = 0;
        memory[ 2213] = 1;
        memory[ 2214] = 1;
        memory[ 2215] = 0;
        memory[ 2216] = 0;
        memory[ 2217] = 0;
        memory[ 2218] = 0;
        memory[ 2219] = 0;
        memory[ 2220] = 0;
        memory[ 2221] = 0;
        memory[ 2222] = 0;
        memory[ 2223] = 0;
        memory[ 2224] = 0;
        memory[ 2225] = 0;
        memory[ 2226] = 1;
        memory[ 2227] = 0;
        memory[ 2228] = 0;
        memory[ 2229] = 0;
        memory[ 2230] = 0;
        memory[ 2231] = 0;
        memory[ 2232] = 1;
        memory[ 2233] = 1;
        memory[ 2234] = 0;
        memory[ 2235] = 0;
        memory[ 2236] = 0;
        memory[ 2237] = 0;
        memory[ 2238] = 0;
        memory[ 2239] = 0;
        memory[ 2240] = 0;
        memory[ 2241] = 0;
        memory[ 2242] = 0;
        memory[ 2243] = 0;
        memory[ 2244] = 0;
        memory[ 2245] = 0;
        memory[ 2246] = 0;
        memory[ 2247] = 1;
        memory[ 2248] = 1;
        memory[ 2249] = 0;
        memory[ 2250] = 0;
        memory[ 2251] = 0;
        memory[ 2252] = 0;
        memory[ 2253] = 0;
        memory[ 2254] = 0;
        memory[ 2255] = 0;
        memory[ 2256] = 1;
        memory[ 2257] = 0;
        memory[ 2258] = 0;
        memory[ 2259] = 0;
        memory[ 2260] = 0;
        memory[ 2261] = 0;
        memory[ 2262] = 0;
        memory[ 2263] = 0;
        memory[ 2264] = 0;
        memory[ 2265] = 0;
        memory[ 2266] = 0;
        memory[ 2267] = 0;
        memory[ 2268] = 1;
        memory[ 2269] = 0;
        memory[ 2270] = 0;
        memory[ 2271] = 0;
        memory[ 2272] = 0;
        memory[ 2273] = 0;
        memory[ 2274] = 0;
        memory[ 2275] = 0;
        memory[ 2276] = 0;
        memory[ 2277] = 0;
        memory[ 2278] = 0;
        memory[ 2279] = 0;
        memory[ 2280] = 0;
        memory[ 2281] = 0;
        memory[ 2282] = 0;
        memory[ 2283] = 0;
        memory[ 2284] = 0;
        memory[ 2285] = 1;
        memory[ 2286] = 1;
        memory[ 2287] = 0;
        memory[ 2288] = 1;
        memory[ 2289] = 0;
        memory[ 2290] = 0;
        memory[ 2291] = 0;
        memory[ 2292] = 0;
        memory[ 2293] = 1;
        memory[ 2294] = 1;
        memory[ 2295] = 0;
        memory[ 2296] = 0;
        memory[ 2297] = 0;
        memory[ 2298] = 0;
        memory[ 2299] = 0;
        memory[ 2300] = 1;
        memory[ 2301] = 1;
        memory[ 2302] = 1;
        memory[ 2303] = 0;
        memory[ 2304] = 0;
        memory[ 2305] = 0;
        memory[ 2306] = 0;
        memory[ 2307] = 0;
        memory[ 2308] = 0;
        memory[ 2309] = 0;
        memory[ 2310] = 0;
        memory[ 2311] = 0;
        memory[ 2312] = 0;
        memory[ 2313] = 0;
        memory[ 2314] = 0;
        memory[ 2315] = 0;
        memory[ 2316] = 0;
        memory[ 2317] = 0;
        memory[ 2318] = 0;
        memory[ 2319] = 0;
        memory[ 2320] = 0;
        memory[ 2321] = 0;
        memory[ 2322] = 0;
        memory[ 2323] = 0;
        memory[ 2324] = 0;
        memory[ 2325] = 0;
        memory[ 2326] = 0;
        memory[ 2327] = 0;
        memory[ 2328] = 0;
        memory[ 2329] = 0;
        memory[ 2330] = 0;
        memory[ 2331] = 0;
        memory[ 2332] = 0;
        memory[ 2333] = 0;
        memory[ 2334] = 0;
        memory[ 2335] = 1;
        memory[ 2336] = 0;
        memory[ 2337] = 0;
        memory[ 2338] = 0;
        memory[ 2339] = 0;
        memory[ 2340] = 1;
        memory[ 2341] = 1;
        memory[ 2342] = 0;
        memory[ 2343] = 1;
        memory[ 2344] = 1;
        memory[ 2345] = 1;
        memory[ 2346] = 1;
        memory[ 2347] = 0;
        memory[ 2348] = 0;
        memory[ 2349] = 0;
        memory[ 2350] = 0;
        memory[ 2351] = 0;
        memory[ 2352] = 0;
        memory[ 2353] = 0;
        memory[ 2354] = 0;
        memory[ 2355] = 0;
        memory[ 2356] = 0;
        memory[ 2357] = 0;
        memory[ 2358] = 0;
        memory[ 2359] = 0;
        memory[ 2360] = 0;
        memory[ 2361] = 0;
        memory[ 2362] = 0;
        memory[ 2363] = 0;
        memory[ 2364] = 0;
        memory[ 2365] = 0;
        memory[ 2366] = 0;
        memory[ 2367] = 0;
        memory[ 2368] = 0;
        memory[ 2369] = 0;
        memory[ 2370] = 0;
        memory[ 2371] = 0;
        memory[ 2372] = 0;
        memory[ 2373] = 0;
        memory[ 2374] = 0;
        memory[ 2375] = 0;
        memory[ 2376] = 0;
        memory[ 2377] = 0;
        memory[ 2378] = 0;
        memory[ 2379] = 0;
        memory[ 2380] = 0;
        memory[ 2381] = 0;
        memory[ 2382] = 1;
        memory[ 2383] = 0;
        memory[ 2384] = 0;
        memory[ 2385] = 0;
        memory[ 2386] = 0;
        memory[ 2387] = 1;
        memory[ 2388] = 0;
        memory[ 2389] = 0;
        memory[ 2390] = 0;
        memory[ 2391] = 0;
        memory[ 2392] = 0;
        memory[ 2393] = 0;
        memory[ 2394] = 0;
        memory[ 2395] = 0;
        memory[ 2396] = 0;
        memory[ 2397] = 0;
        memory[ 2398] = 0;
        memory[ 2399] = 0;
        memory[ 2400] = 0;
        memory[ 2401] = 1;
        memory[ 2402] = 1;
        memory[ 2403] = 0;
        memory[ 2404] = 0;
        memory[ 2405] = 0;
        memory[ 2406] = 0;
        memory[ 2407] = 0;
        memory[ 2408] = 0;
        memory[ 2409] = 0;
        memory[ 2410] = 0;
        memory[ 2411] = 0;
        memory[ 2412] = 0;
        memory[ 2413] = 0;
        memory[ 2414] = 0;
        memory[ 2415] = 0;
        memory[ 2416] = 0;
        memory[ 2417] = 1;
        memory[ 2418] = 0;
        memory[ 2419] = 1;
        memory[ 2420] = 0;
        memory[ 2421] = 0;
        memory[ 2422] = 0;
        memory[ 2423] = 0;
        memory[ 2424] = 0;
        memory[ 2425] = 0;
        memory[ 2426] = 0;
        memory[ 2427] = 0;
        memory[ 2428] = 0;
        memory[ 2429] = 0;
        memory[ 2430] = 0;
        memory[ 2431] = 0;
        memory[ 2432] = 0;
        memory[ 2433] = 0;
        memory[ 2434] = 0;
        memory[ 2435] = 0;
        memory[ 2436] = 0;
        memory[ 2437] = 0;
        memory[ 2438] = 0;
        memory[ 2439] = 0;
        memory[ 2440] = 0;
        memory[ 2441] = 0;
        memory[ 2442] = 0;
        memory[ 2443] = 0;
        memory[ 2444] = 0;
        memory[ 2445] = 0;
        memory[ 2446] = 0;
        memory[ 2447] = 0;
        memory[ 2448] = 0;
        memory[ 2449] = 0;
        memory[ 2450] = 0;
        memory[ 2451] = 0;
        memory[ 2452] = 0;
        memory[ 2453] = 0;
        memory[ 2454] = 0;
        memory[ 2455] = 0;
        memory[ 2456] = 0;
        memory[ 2457] = 0;
        memory[ 2458] = 0;
        memory[ 2459] = 0;
        memory[ 2460] = 1;
        memory[ 2461] = 0;
        memory[ 2462] = 0;
        memory[ 2463] = 0;
        memory[ 2464] = 0;
        memory[ 2465] = 0;
        memory[ 2466] = 0;
        memory[ 2467] = 0;
        memory[ 2468] = 0;
        memory[ 2469] = 0;
        memory[ 2470] = 1;
        memory[ 2471] = 0;
        memory[ 2472] = 0;
        memory[ 2473] = 1;
        memory[ 2474] = 0;
        memory[ 2475] = 0;
        memory[ 2476] = 0;
        memory[ 2477] = 0;
        memory[ 2478] = 0;
        memory[ 2479] = 1;
        memory[ 2480] = 0;
        memory[ 2481] = 0;
        memory[ 2482] = 1;
        memory[ 2483] = 0;
        memory[ 2484] = 0;
        memory[ 2485] = 0;
        memory[ 2486] = 0;
        memory[ 2487] = 0;
        memory[ 2488] = 0;
        memory[ 2489] = 0;
        memory[ 2490] = 0;
        memory[ 2491] = 0;
        memory[ 2492] = 0;
        memory[ 2493] = 0;
        memory[ 2494] = 1;
        memory[ 2495] = 0;
        memory[ 2496] = 0;
        memory[ 2497] = 0;
        memory[ 2498] = 0;
        memory[ 2499] = 0;
        memory[ 2500] = 0;
        memory[ 2501] = 0;
        memory[ 2502] = 0;
        memory[ 2503] = 0;
        memory[ 2504] = 0;
        memory[ 2505] = 0;
        memory[ 2506] = 0;
        memory[ 2507] = 0;
        memory[ 2508] = 0;
        memory[ 2509] = 0;
        memory[ 2510] = 0;
        memory[ 2511] = 0;
        memory[ 2512] = 0;
        memory[ 2513] = 0;
        memory[ 2514] = 1;
        memory[ 2515] = 0;
        memory[ 2516] = 0;
        memory[ 2517] = 0;
        memory[ 2518] = 0;
        memory[ 2519] = 0;
        memory[ 2520] = 0;
        memory[ 2521] = 0;
        memory[ 2522] = 0;
        memory[ 2523] = 0;
        memory[ 2524] = 0;
        memory[ 2525] = 0;
        memory[ 2526] = 0;
        memory[ 2527] = 0;
        memory[ 2528] = 1;
        memory[ 2529] = 1;
        memory[ 2530] = 0;
        memory[ 2531] = 0;
        memory[ 2532] = 0;
        memory[ 2533] = 0;
        memory[ 2534] = 0;
        memory[ 2535] = 0;
        memory[ 2536] = 0;
        memory[ 2537] = 0;
        memory[ 2538] = 0;
        memory[ 2539] = 0;
        memory[ 2540] = 0;
        memory[ 2541] = 0;
        memory[ 2542] = 0;
        memory[ 2543] = 0;
        memory[ 2544] = 0;
        memory[ 2545] = 0;
        memory[ 2546] = 0;
        memory[ 2547] = 0;
        memory[ 2548] = 0;
        memory[ 2549] = 0;
        memory[ 2550] = 0;
        memory[ 2551] = 0;
        memory[ 2552] = 0;
        memory[ 2553] = 0;
        memory[ 2554] = 0;
        memory[ 2555] = 0;
        memory[ 2556] = 0;
        memory[ 2557] = 0;
        memory[ 2558] = 0;
        memory[ 2559] = 0;
        memory[ 2560] = 0;
        memory[ 2561] = 0;
        memory[ 2562] = 0;
        memory[ 2563] = 0;
        memory[ 2564] = 0;
        memory[ 2565] = 0;
        memory[ 2566] = 0;
        memory[ 2567] = 0;
        memory[ 2568] = 0;
        memory[ 2569] = 0;
        memory[ 2570] = 1;
        memory[ 2571] = 0;
        memory[ 2572] = 0;
        memory[ 2573] = 0;
        memory[ 2574] = 0;
        memory[ 2575] = 0;
        memory[ 2576] = 0;
        memory[ 2577] = 0;
        memory[ 2578] = 0;
        memory[ 2579] = 0;
        memory[ 2580] = 0;
        memory[ 2581] = 0;
        memory[ 2582] = 0;
        memory[ 2583] = 0;
        memory[ 2584] = 0;
        memory[ 2585] = 0;
        memory[ 2586] = 0;
        memory[ 2587] = 0;
        memory[ 2588] = 0;
        memory[ 2589] = 0;
        memory[ 2590] = 0;
        memory[ 2591] = 0;
        memory[ 2592] = 1;
        memory[ 2593] = 0;
        memory[ 2594] = 1;
        memory[ 2595] = 0;
        memory[ 2596] = 0;
        memory[ 2597] = 0;
        memory[ 2598] = 0;
        memory[ 2599] = 0;
        memory[ 2600] = 0;
        memory[ 2601] = 0;
        memory[ 2602] = 0;
        memory[ 2603] = 0;
        memory[ 2604] = 0;
        memory[ 2605] = 0;
        memory[ 2606] = 0;
        memory[ 2607] = 0;
        memory[ 2608] = 1;
        memory[ 2609] = 1;
        memory[ 2610] = 1;
        memory[ 2611] = 1;
        memory[ 2612] = 1;
        memory[ 2613] = 0;
        memory[ 2614] = 0;
        memory[ 2615] = 0;
        memory[ 2616] = 0;
        memory[ 2617] = 0;
        memory[ 2618] = 0;
        memory[ 2619] = 0;
        memory[ 2620] = 0;
        memory[ 2621] = 0;
        memory[ 2622] = 0;
        memory[ 2623] = 0;
        memory[ 2624] = 0;
        memory[ 2625] = 0;
        memory[ 2626] = 0;
        memory[ 2627] = 0;
        memory[ 2628] = 0;
        memory[ 2629] = 0;
        memory[ 2630] = 0;
        memory[ 2631] = 0;
        memory[ 2632] = 0;
        memory[ 2633] = 0;
        memory[ 2634] = 0;
        memory[ 2635] = 0;
        memory[ 2636] = 0;
        memory[ 2637] = 0;
        memory[ 2638] = 0;
        memory[ 2639] = 0;
        memory[ 2640] = 0;
        memory[ 2641] = 0;
        memory[ 2642] = 0;
        memory[ 2643] = 0;
        memory[ 2644] = 0;
        memory[ 2645] = 0;
        memory[ 2646] = 0;
        memory[ 2647] = 0;
        memory[ 2648] = 0;
        memory[ 2649] = 0;
        memory[ 2650] = 0;
        memory[ 2651] = 1;
        memory[ 2652] = 0;
        memory[ 2653] = 0;
        memory[ 2654] = 0;
        memory[ 2655] = 0;
        memory[ 2656] = 0;
        memory[ 2657] = 0;
        memory[ 2658] = 0;
        memory[ 2659] = 0;
        memory[ 2660] = 0;
        memory[ 2661] = 0;
        memory[ 2662] = 0;
        memory[ 2663] = 0;
        memory[ 2664] = 0;
        memory[ 2665] = 0;
        memory[ 2666] = 0;
        memory[ 2667] = 0;
        memory[ 2668] = 0;
        memory[ 2669] = 0;
        memory[ 2670] = 0;
        memory[ 2671] = 0;
        memory[ 2672] = 0;
        memory[ 2673] = 0;
        memory[ 2674] = 0;
        memory[ 2675] = 0;
        memory[ 2676] = 0;
        memory[ 2677] = 0;
        memory[ 2678] = 0;
        memory[ 2679] = 0;
        memory[ 2680] = 0;
        memory[ 2681] = 0;
        memory[ 2682] = 0;
        memory[ 2683] = 0;
        memory[ 2684] = 0;
        memory[ 2685] = 0;
        memory[ 2686] = 0;
        memory[ 2687] = 0;
        memory[ 2688] = 0;
        memory[ 2689] = 0;
        memory[ 2690] = 0;
        memory[ 2691] = 1;
        memory[ 2692] = 0;
        memory[ 2693] = 0;
        memory[ 2694] = 0;
        memory[ 2695] = 0;
        memory[ 2696] = 0;
        memory[ 2697] = 0;
        memory[ 2698] = 0;
        memory[ 2699] = 0;
        memory[ 2700] = 1;
        memory[ 2701] = 0;
        memory[ 2702] = 1;
        memory[ 2703] = 0;
        memory[ 2704] = 0;
        memory[ 2705] = 0;
        memory[ 2706] = 0;
        memory[ 2707] = 0;
        memory[ 2708] = 1;
        memory[ 2709] = 0;
        memory[ 2710] = 0;
        memory[ 2711] = 0;
        memory[ 2712] = 0;
        memory[ 2713] = 0;
        memory[ 2714] = 0;
        memory[ 2715] = 0;
        memory[ 2716] = 0;
        memory[ 2717] = 0;
        memory[ 2718] = 0;
        memory[ 2719] = 1;
        memory[ 2720] = 0;
        memory[ 2721] = 0;
        memory[ 2722] = 0;
        memory[ 2723] = 0;
        memory[ 2724] = 0;
        memory[ 2725] = 0;
        memory[ 2726] = 0;
        memory[ 2727] = 0;
        memory[ 2728] = 0;
        memory[ 2729] = 0;
        memory[ 2730] = 0;
        memory[ 2731] = 0;
        memory[ 2732] = 0;
        memory[ 2733] = 0;
        memory[ 2734] = 0;
        memory[ 2735] = 0;
        memory[ 2736] = 0;
        memory[ 2737] = 0;
        memory[ 2738] = 0;
        memory[ 2739] = 0;
        memory[ 2740] = 0;
        memory[ 2741] = 0;
        memory[ 2742] = 0;
        memory[ 2743] = 0;
        memory[ 2744] = 0;
        memory[ 2745] = 0;
        memory[ 2746] = 0;
        memory[ 2747] = 0;
        memory[ 2748] = 0;
        memory[ 2749] = 0;
        memory[ 2750] = 0;
        memory[ 2751] = 0;
        memory[ 2752] = 0;
        memory[ 2753] = 0;
        memory[ 2754] = 0;
        memory[ 2755] = 0;
        memory[ 2756] = 0;
        memory[ 2757] = 0;
        memory[ 2758] = 0;
        memory[ 2759] = 0;
        memory[ 2760] = 0;
        memory[ 2761] = 0;
        memory[ 2762] = 0;
        memory[ 2763] = 0;
        memory[ 2764] = 0;
        memory[ 2765] = 0;
        memory[ 2766] = 0;
        memory[ 2767] = 0;
        memory[ 2768] = 0;
        memory[ 2769] = 0;
        memory[ 2770] = 0;
        memory[ 2771] = 0;
        memory[ 2772] = 0;
        memory[ 2773] = 0;
        memory[ 2774] = 1;
        memory[ 2775] = 0;
        memory[ 2776] = 0;
        memory[ 2777] = 1;
        memory[ 2778] = 0;
        memory[ 2779] = 0;
        memory[ 2780] = 0;
        memory[ 2781] = 0;
        memory[ 2782] = 0;
        memory[ 2783] = 0;
        memory[ 2784] = 0;
        memory[ 2785] = 0;
        memory[ 2786] = 0;
        memory[ 2787] = 0;
        memory[ 2788] = 0;
        memory[ 2789] = 0;
        memory[ 2790] = 0;
        memory[ 2791] = 0;
        memory[ 2792] = 0;
        memory[ 2793] = 0;
        memory[ 2794] = 0;
        memory[ 2795] = 0;
        memory[ 2796] = 0;
        memory[ 2797] = 1;
        memory[ 2798] = 0;
        memory[ 2799] = 0;
        memory[ 2800] = 1;
        memory[ 2801] = 0;
        memory[ 2802] = 0;
        memory[ 2803] = 0;
        memory[ 2804] = 0;
        memory[ 2805] = 0;
        memory[ 2806] = 0;
        memory[ 2807] = 0;
        memory[ 2808] = 0;
        memory[ 2809] = 0;
        memory[ 2810] = 0;
        memory[ 2811] = 0;
        memory[ 2812] = 0;
        memory[ 2813] = 0;
        memory[ 2814] = 0;
        memory[ 2815] = 0;
        memory[ 2816] = 0;
        memory[ 2817] = 0;
        memory[ 2818] = 0;
        memory[ 2819] = 1;
        memory[ 2820] = 0;
        memory[ 2821] = 0;
        memory[ 2822] = 0;
        memory[ 2823] = 0;
        memory[ 2824] = 0;
        memory[ 2825] = 0;
        memory[ 2826] = 0;
        memory[ 2827] = 0;
        memory[ 2828] = 0;
        memory[ 2829] = 0;
        memory[ 2830] = 0;
        memory[ 2831] = 0;
        memory[ 2832] = 0;
        memory[ 2833] = 0;
        memory[ 2834] = 0;
        memory[ 2835] = 0;
        memory[ 2836] = 0;
        memory[ 2837] = 0;
        memory[ 2838] = 0;
        memory[ 2839] = 0;
        memory[ 2840] = 0;
        memory[ 2841] = 0;
        memory[ 2842] = 0;
        memory[ 2843] = 0;
        memory[ 2844] = 0;
        memory[ 2845] = 0;
        memory[ 2846] = 0;
        memory[ 2847] = 0;
        memory[ 2848] = 0;
        memory[ 2849] = 0;
        memory[ 2850] = 0;
        memory[ 2851] = 0;
        memory[ 2852] = 0;
        memory[ 2853] = 0;
        memory[ 2854] = 0;
        memory[ 2855] = 0;
        memory[ 2856] = 0;
        memory[ 2857] = 0;
        memory[ 2858] = 0;
        memory[ 2859] = 0;
        memory[ 2860] = 0;
        memory[ 2861] = 0;
        memory[ 2862] = 0;
        memory[ 2863] = 0;
        memory[ 2864] = 0;
        memory[ 2865] = 0;
        memory[ 2866] = 0;
        memory[ 2867] = 0;
        memory[ 2868] = 1;
        memory[ 2869] = 0;
        memory[ 2870] = 0;
        memory[ 2871] = 0;
        memory[ 2872] = 0;
        memory[ 2873] = 0;
        memory[ 2874] = 0;
        memory[ 2875] = 0;
        memory[ 2876] = 1;
        memory[ 2877] = 0;
        memory[ 2878] = 1;
        memory[ 2879] = 0;
        memory[ 2880] = 0;
        memory[ 2881] = 0;
        memory[ 2882] = 0;
        memory[ 2883] = 0;
        memory[ 2884] = 0;
        memory[ 2885] = 0;
        memory[ 2886] = 0;
        memory[ 2887] = 0;
        memory[ 2888] = 0;
        memory[ 2889] = 1;
        memory[ 2890] = 0;
        memory[ 2891] = 0;
        memory[ 2892] = 0;
        memory[ 2893] = 0;
        memory[ 2894] = 0;
        memory[ 2895] = 0;
        memory[ 2896] = 0;
        memory[ 2897] = 0;
        memory[ 2898] = 0;
        memory[ 2899] = 0;
        memory[ 2900] = 0;
        memory[ 2901] = 0;
        memory[ 2902] = 0;
        memory[ 2903] = 0;
        memory[ 2904] = 0;
        memory[ 2905] = 0;
        memory[ 2906] = 0;
        memory[ 2907] = 0;
        memory[ 2908] = 0;
        memory[ 2909] = 0;
        memory[ 2910] = 0;
        memory[ 2911] = 0;
        memory[ 2912] = 0;
        memory[ 2913] = 0;
        memory[ 2914] = 0;
        memory[ 2915] = 0;
        memory[ 2916] = 0;
        memory[ 2917] = 0;
        memory[ 2918] = 0;
        memory[ 2919] = 0;
        memory[ 2920] = 0;
        memory[ 2921] = 0;
        memory[ 2922] = 0;
        memory[ 2923] = 0;
        memory[ 2924] = 0;
        memory[ 2925] = 0;
        memory[ 2926] = 0;
        memory[ 2927] = 0;
        memory[ 2928] = 0;
        memory[ 2929] = 0;
        memory[ 2930] = 0;
        memory[ 2931] = 0;
        memory[ 2932] = 0;
        memory[ 2933] = 0;
        memory[ 2934] = 1;
        memory[ 2935] = 0;
        memory[ 2936] = 0;
        memory[ 2937] = 0;
        memory[ 2938] = 0;
        memory[ 2939] = 0;
        memory[ 2940] = 0;
        memory[ 2941] = 0;
        memory[ 2942] = 0;
        memory[ 2943] = 0;
        memory[ 2944] = 0;
        memory[ 2945] = 0;
        memory[ 2946] = 0;
        memory[ 2947] = 0;
        memory[ 2948] = 0;
        memory[ 2949] = 0;
        memory[ 2950] = 0;
        memory[ 2951] = 0;
        memory[ 2952] = 0;
        memory[ 2953] = 0;
        memory[ 2954] = 0;
        memory[ 2955] = 0;
        memory[ 2956] = 1;
        memory[ 2957] = 1;
        memory[ 2958] = 0;
        memory[ 2959] = 0;
        memory[ 2960] = 0;
        memory[ 2961] = 0;
        memory[ 2962] = 0;
        memory[ 2963] = 1;
        memory[ 2964] = 1;
        memory[ 2965] = 0;
        memory[ 2966] = 0;
        memory[ 2967] = 0;
        memory[ 2968] = 0;
        memory[ 2969] = 0;
        memory[ 2970] = 0;
        memory[ 2971] = 0;
        memory[ 2972] = 0;
        memory[ 2973] = 0;
        memory[ 2974] = 0;
        memory[ 2975] = 0;
        memory[ 2976] = 0;
        memory[ 2977] = 1;
        memory[ 2978] = 0;
        memory[ 2979] = 0;
        memory[ 2980] = 1;
        memory[ 2981] = 0;
        memory[ 2982] = 0;
        memory[ 2983] = 0;
        memory[ 2984] = 0;
        memory[ 2985] = 0;
        memory[ 2986] = 0;
        memory[ 2987] = 0;
        memory[ 2988] = 0;
        memory[ 2989] = 0;
        memory[ 2990] = 0;
        memory[ 2991] = 0;
        memory[ 2992] = 0;
        memory[ 2993] = 0;
        memory[ 2994] = 0;
        memory[ 2995] = 0;
        memory[ 2996] = 0;
        memory[ 2997] = 0;
        memory[ 2998] = 0;
        memory[ 2999] = 0;
        memory[ 3000] = 0;
        memory[ 3001] = 0;
        memory[ 3002] = 0;
        memory[ 3003] = 0;
        memory[ 3004] = 0;
        memory[ 3005] = 0;
        memory[ 3006] = 0;
        memory[ 3007] = 0;
        memory[ 3008] = 0;
        memory[ 3009] = 0;
        memory[ 3010] = 0;
        memory[ 3011] = 1;
        memory[ 3012] = 1;
        memory[ 3013] = 0;
        memory[ 3014] = 0;
        memory[ 3015] = 0;
        memory[ 3016] = 0;
        memory[ 3017] = 0;
        memory[ 3018] = 0;
        memory[ 3019] = 0;
        memory[ 3020] = 0;
        memory[ 3021] = 1;
        memory[ 3022] = 0;
        memory[ 3023] = 0;
        memory[ 3024] = 0;
        memory[ 3025] = 0;
        memory[ 3026] = 0;
        memory[ 3027] = 0;
        memory[ 3028] = 0;
        memory[ 3029] = 0;
        memory[ 3030] = 0;
        memory[ 3031] = 0;
        memory[ 3032] = 0;
        memory[ 3033] = 0;
        memory[ 3034] = 0;
        memory[ 3035] = 0;
        memory[ 3036] = 0;
        memory[ 3037] = 0;
        memory[ 3038] = 0;
        memory[ 3039] = 0;
        memory[ 3040] = 0;
        memory[ 3041] = 1;
        memory[ 3042] = 0;
        memory[ 3043] = 0;
        memory[ 3044] = 1;
        memory[ 3045] = 1;
        memory[ 3046] = 0;
        memory[ 3047] = 0;
        memory[ 3048] = 1;
        memory[ 3049] = 0;
        memory[ 3050] = 0;
        memory[ 3051] = 0;
        memory[ 3052] = 0;
        memory[ 3053] = 0;
        memory[ 3054] = 0;
        memory[ 3055] = 0;
        memory[ 3056] = 0;
        memory[ 3057] = 0;
        memory[ 3058] = 0;
        memory[ 3059] = 0;
        memory[ 3060] = 1;
        memory[ 3061] = 0;
        memory[ 3062] = 0;
        memory[ 3063] = 0;
        memory[ 3064] = 0;
        memory[ 3065] = 0;
        memory[ 3066] = 0;
        memory[ 3067] = 0;
        memory[ 3068] = 0;
        memory[ 3069] = 0;
        memory[ 3070] = 1;
        memory[ 3071] = 0;
        memory[ 3072] = 0;
        memory[ 3073] = 0;
        memory[ 3074] = 0;
        memory[ 3075] = 0;
        memory[ 3076] = 0;
        memory[ 3077] = 0;
        memory[ 3078] = 0;
        memory[ 3079] = 0;
        memory[ 3080] = 0;
        memory[ 3081] = 0;
        memory[ 3082] = 0;
        memory[ 3083] = 0;
        memory[ 3084] = 0;
        memory[ 3085] = 0;
        memory[ 3086] = 0;
        memory[ 3087] = 0;
        memory[ 3088] = 0;
        memory[ 3089] = 0;
        memory[ 3090] = 0;
        memory[ 3091] = 1;
        memory[ 3092] = 0;
        memory[ 3093] = 0;
        memory[ 3094] = 0;
        memory[ 3095] = 0;
        memory[ 3096] = 0;
        memory[ 3097] = 0;
        memory[ 3098] = 0;
        memory[ 3099] = 0;
        memory[ 3100] = 0;
        memory[ 3101] = 0;
        memory[ 3102] = 0;
        memory[ 3103] = 0;
        memory[ 3104] = 0;
        memory[ 3105] = 0;
        memory[ 3106] = 0;
        memory[ 3107] = 0;
        memory[ 3108] = 0;
        memory[ 3109] = 0;
        memory[ 3110] = 1;
        memory[ 3111] = 1;
        memory[ 3112] = 0;
        memory[ 3113] = 0;
        memory[ 3114] = 0;
        memory[ 3115] = 0;
        memory[ 3116] = 0;
        memory[ 3117] = 0;
        memory[ 3118] = 0;
        memory[ 3119] = 0;
        memory[ 3120] = 0;
        memory[ 3121] = 0;
        memory[ 3122] = 0;
        memory[ 3123] = 0;
        memory[ 3124] = 0;
        memory[ 3125] = 0;
        memory[ 3126] = 0;
        memory[ 3127] = 0;
        memory[ 3128] = 0;
        memory[ 3129] = 0;
        memory[ 3130] = 0;
        memory[ 3131] = 0;
        memory[ 3132] = 0;
        memory[ 3133] = 0;
        memory[ 3134] = 0;
        memory[ 3135] = 1;
        memory[ 3136] = 1;
        memory[ 3137] = 1;
        memory[ 3138] = 1;
        memory[ 3139] = 0;
        memory[ 3140] = 1;
        memory[ 3141] = 0;
        memory[ 3142] = 0;
        memory[ 3143] = 0;
        memory[ 3144] = 0;
        memory[ 3145] = 0;
        memory[ 3146] = 0;
        memory[ 3147] = 0;
        memory[ 3148] = 0;
        memory[ 3149] = 0;
        memory[ 3150] = 0;
        memory[ 3151] = 0;
        memory[ 3152] = 0;
        memory[ 3153] = 0;
        memory[ 3154] = 0;
        memory[ 3155] = 0;
        memory[ 3156] = 0;
        memory[ 3157] = 0;
        memory[ 3158] = 0;
        memory[ 3159] = 0;
        memory[ 3160] = 1;
        memory[ 3161] = 0;
        memory[ 3162] = 0;
        memory[ 3163] = 0;
        memory[ 3164] = 0;
        memory[ 3165] = 0;
        memory[ 3166] = 0;
        memory[ 3167] = 0;
        memory[ 3168] = 0;
        memory[ 3169] = 0;
        memory[ 3170] = 0;
        memory[ 3171] = 0;
        memory[ 3172] = 0;
        memory[ 3173] = 1;
        memory[ 3174] = 0;
        memory[ 3175] = 0;
        memory[ 3176] = 0;
        memory[ 3177] = 0;
        memory[ 3178] = 0;
        memory[ 3179] = 1;
        memory[ 3180] = 0;
        memory[ 3181] = 0;
        memory[ 3182] = 0;
        memory[ 3183] = 0;
        memory[ 3184] = 1;
        memory[ 3185] = 1;
        memory[ 3186] = 0;
        memory[ 3187] = 0;
        memory[ 3188] = 1;
        memory[ 3189] = 0;
        memory[ 3190] = 0;
        memory[ 3191] = 0;
        memory[ 3192] = 1;
        memory[ 3193] = 0;
        memory[ 3194] = 0;
        memory[ 3195] = 0;
        memory[ 3196] = 0;
        memory[ 3197] = 0;
        memory[ 3198] = 0;
        memory[ 3199] = 0;
        memory[ 3200] = 0;
        memory[ 3201] = 0;
        memory[ 3202] = 0;
        memory[ 3203] = 0;
        memory[ 3204] = 0;
        memory[ 3205] = 0;
        memory[ 3206] = 0;
        memory[ 3207] = 0;
        memory[ 3208] = 0;
        memory[ 3209] = 0;
        memory[ 3210] = 0;
        memory[ 3211] = 0;
        memory[ 3212] = 0;
        memory[ 3213] = 0;
        memory[ 3214] = 0;
        memory[ 3215] = 0;
        memory[ 3216] = 0;
        memory[ 3217] = 0;
        memory[ 3218] = 0;
        memory[ 3219] = 0;
        memory[ 3220] = 0;
        memory[ 3221] = 0;
        memory[ 3222] = 0;
        memory[ 3223] = 0;
        memory[ 3224] = 0;
        memory[ 3225] = 0;
        memory[ 3226] = 0;
        memory[ 3227] = 0;
        memory[ 3228] = 0;
        memory[ 3229] = 1;
        memory[ 3230] = 0;
        memory[ 3231] = 1;
        memory[ 3232] = 0;
        memory[ 3233] = 0;
        memory[ 3234] = 0;
        memory[ 3235] = 0;
        memory[ 3236] = 0;
        memory[ 3237] = 0;
        memory[ 3238] = 0;
        memory[ 3239] = 0;
        memory[ 3240] = 0;
        memory[ 3241] = 0;
        memory[ 3242] = 0;
        memory[ 3243] = 0;
        memory[ 3244] = 0;
        memory[ 3245] = 0;
        memory[ 3246] = 0;
        memory[ 3247] = 0;
        memory[ 3248] = 0;
        memory[ 3249] = 0;
        memory[ 3250] = 0;
        memory[ 3251] = 0;
        memory[ 3252] = 1;
        memory[ 3253] = 0;
        memory[ 3254] = 0;
        memory[ 3255] = 0;
        memory[ 3256] = 0;
        memory[ 3257] = 0;
        memory[ 3258] = 0;
        memory[ 3259] = 0;
        memory[ 3260] = 0;
        memory[ 3261] = 0;
        memory[ 3262] = 0;
        memory[ 3263] = 0;
        memory[ 3264] = 0;
        memory[ 3265] = 0;
        memory[ 3266] = 0;
        memory[ 3267] = 1;
        memory[ 3268] = 0;
        memory[ 3269] = 0;
        memory[ 3270] = 0;
        memory[ 3271] = 0;
        memory[ 3272] = 0;
        memory[ 3273] = 0;
        memory[ 3274] = 1;
        memory[ 3275] = 1;
        memory[ 3276] = 0;
        memory[ 3277] = 0;
        memory[ 3278] = 0;
        memory[ 3279] = 0;
        memory[ 3280] = 0;
        memory[ 3281] = 0;
        memory[ 3282] = 0;
        memory[ 3283] = 1;
        memory[ 3284] = 0;
        memory[ 3285] = 0;
        memory[ 3286] = 0;
        memory[ 3287] = 0;
        memory[ 3288] = 0;
        memory[ 3289] = 0;
        memory[ 3290] = 0;
        memory[ 3291] = 0;
        memory[ 3292] = 0;
        memory[ 3293] = 0;
        memory[ 3294] = 0;
        memory[ 3295] = 0;
        memory[ 3296] = 0;
        memory[ 3297] = 0;
        memory[ 3298] = 0;
        memory[ 3299] = 0;
        memory[ 3300] = 0;
        memory[ 3301] = 0;
        memory[ 3302] = 0;
        memory[ 3303] = 0;
        memory[ 3304] = 0;
        memory[ 3305] = 0;
        memory[ 3306] = 0;
        memory[ 3307] = 0;
        memory[ 3308] = 0;
        memory[ 3309] = 1;
        memory[ 3310] = 1;
        memory[ 3311] = 1;
        memory[ 3312] = 0;
        memory[ 3313] = 0;
        memory[ 3314] = 0;
        memory[ 3315] = 0;
        memory[ 3316] = 0;
        memory[ 3317] = 0;
        memory[ 3318] = 0;
        memory[ 3319] = 0;
        memory[ 3320] = 0;
        memory[ 3321] = 0;
        memory[ 3322] = 0;
        memory[ 3323] = 0;
        memory[ 3324] = 0;
        memory[ 3325] = 0;
        memory[ 3326] = 0;
        memory[ 3327] = 0;
        memory[ 3328] = 0;
        memory[ 3329] = 0;
        memory[ 3330] = 0;
        memory[ 3331] = 0;
        memory[ 3332] = 0;
        memory[ 3333] = 1;
        memory[ 3334] = 0;
        memory[ 3335] = 0;
        memory[ 3336] = 0;
        memory[ 3337] = 0;
        memory[ 3338] = 0;
        memory[ 3339] = 1;
        memory[ 3340] = 1;
        memory[ 3341] = 0;
        memory[ 3342] = 0;
        memory[ 3343] = 0;
        memory[ 3344] = 0;
        memory[ 3345] = 0;
        memory[ 3346] = 0;
        memory[ 3347] = 0;
        memory[ 3348] = 0;
        memory[ 3349] = 0;
        memory[ 3350] = 0;
        memory[ 3351] = 0;
        memory[ 3352] = 1;
        memory[ 3353] = 0;
        memory[ 3354] = 0;
        memory[ 3355] = 0;
        memory[ 3356] = 0;
        memory[ 3357] = 0;
        memory[ 3358] = 0;
        memory[ 3359] = 0;
        memory[ 3360] = 0;
        memory[ 3361] = 1;
        memory[ 3362] = 0;
        memory[ 3363] = 0;
        memory[ 3364] = 1;
        memory[ 3365] = 0;
        memory[ 3366] = 0;
        memory[ 3367] = 0;
        memory[ 3368] = 0;
        memory[ 3369] = 0;
        memory[ 3370] = 1;
        memory[ 3371] = 0;
        memory[ 3372] = 0;
        memory[ 3373] = 0;
        memory[ 3374] = 0;
        memory[ 3375] = 0;
        memory[ 3376] = 0;
        memory[ 3377] = 0;
        memory[ 3378] = 0;
        memory[ 3379] = 0;
        memory[ 3380] = 0;
        memory[ 3381] = 0;
        memory[ 3382] = 0;
        memory[ 3383] = 0;
        memory[ 3384] = 0;
        memory[ 3385] = 0;
        memory[ 3386] = 1;
        memory[ 3387] = 0;
        memory[ 3388] = 0;
        memory[ 3389] = 0;
        memory[ 3390] = 0;
        memory[ 3391] = 0;
        memory[ 3392] = 0;
        memory[ 3393] = 0;
        memory[ 3394] = 0;
        memory[ 3395] = 0;
        memory[ 3396] = 0;
        memory[ 3397] = 0;
        memory[ 3398] = 0;
        memory[ 3399] = 0;
        memory[ 3400] = 0;
        memory[ 3401] = 0;
        memory[ 3402] = 1;
        memory[ 3403] = 0;
        memory[ 3404] = 0;
        memory[ 3405] = 0;
        memory[ 3406] = 0;
        memory[ 3407] = 1;
        memory[ 3408] = 0;
        memory[ 3409] = 0;
        memory[ 3410] = 0;
        memory[ 3411] = 0;
        memory[ 3412] = 0;
        memory[ 3413] = 0;
        memory[ 3414] = 1;
        memory[ 3415] = 0;
        memory[ 3416] = 0;
        memory[ 3417] = 0;
        memory[ 3418] = 0;
        memory[ 3419] = 0;
        memory[ 3420] = 0;
        memory[ 3421] = 0;
        memory[ 3422] = 1;
        memory[ 3423] = 0;
        memory[ 3424] = 0;
        memory[ 3425] = 0;
        memory[ 3426] = 0;
        memory[ 3427] = 0;
        memory[ 3428] = 0;
        memory[ 3429] = 0;
        memory[ 3430] = 0;
        memory[ 3431] = 0;
        memory[ 3432] = 0;
        memory[ 3433] = 0;
        memory[ 3434] = 0;
        memory[ 3435] = 0;
        memory[ 3436] = 0;
        memory[ 3437] = 0;
        memory[ 3438] = 1;
        memory[ 3439] = 0;
        memory[ 3440] = 0;
        memory[ 3441] = 0;
        memory[ 3442] = 0;
        memory[ 3443] = 0;
        memory[ 3444] = 0;
        memory[ 3445] = 0;
        memory[ 3446] = 0;
        memory[ 3447] = 0;
        memory[ 3448] = 0;
        memory[ 3449] = 1;
        memory[ 3450] = 0;
        memory[ 3451] = 0;
        memory[ 3452] = 0;
        memory[ 3453] = 0;
        memory[ 3454] = 1;
        memory[ 3455] = 1;
        memory[ 3456] = 0;
        memory[ 3457] = 0;
        memory[ 3458] = 1;
        memory[ 3459] = 1;
        memory[ 3460] = 1;
        memory[ 3461] = 1;
        memory[ 3462] = 0;
        memory[ 3463] = 0;
        memory[ 3464] = 0;
        memory[ 3465] = 0;
        memory[ 3466] = 0;
        memory[ 3467] = 0;
        memory[ 3468] = 0;
        memory[ 3469] = 0;
        memory[ 3470] = 0;
        memory[ 3471] = 0;
        memory[ 3472] = 0;
        memory[ 3473] = 0;
        memory[ 3474] = 0;
        memory[ 3475] = 0;
        memory[ 3476] = 1;
        memory[ 3477] = 0;
        memory[ 3478] = 0;
        memory[ 3479] = 0;
        memory[ 3480] = 0;
        memory[ 3481] = 0;
        memory[ 3482] = 0;
        memory[ 3483] = 0;
        memory[ 3484] = 0;
        memory[ 3485] = 0;
        memory[ 3486] = 0;
        memory[ 3487] = 0;
        memory[ 3488] = 0;
        memory[ 3489] = 0;
        memory[ 3490] = 0;
        memory[ 3491] = 0;
        memory[ 3492] = 0;
        memory[ 3493] = 0;
        memory[ 3494] = 0;
        memory[ 3495] = 0;
        memory[ 3496] = 0;
        memory[ 3497] = 1;
        memory[ 3498] = 1;
        memory[ 3499] = 0;
        memory[ 3500] = 0;
        memory[ 3501] = 0;
        memory[ 3502] = 0;
        memory[ 3503] = 0;
        memory[ 3504] = 0;
        memory[ 3505] = 0;
        memory[ 3506] = 0;
        memory[ 3507] = 0;
        memory[ 3508] = 1;
        memory[ 3509] = 0;
        memory[ 3510] = 0;
        memory[ 3511] = 0;
        memory[ 3512] = 0;
        memory[ 3513] = 1;
        memory[ 3514] = 0;
        memory[ 3515] = 0;
        memory[ 3516] = 0;
        memory[ 3517] = 0;
        memory[ 3518] = 0;
        memory[ 3519] = 0;
        memory[ 3520] = 0;
        memory[ 3521] = 0;
        memory[ 3522] = 0;
        memory[ 3523] = 0;
        memory[ 3524] = 0;
        memory[ 3525] = 0;
        memory[ 3526] = 0;
        memory[ 3527] = 1;
        memory[ 3528] = 0;
        memory[ 3529] = 0;
        memory[ 3530] = 0;
        memory[ 3531] = 0;
        memory[ 3532] = 0;
        memory[ 3533] = 0;
        memory[ 3534] = 0;
        memory[ 3535] = 0;
        memory[ 3536] = 0;
        memory[ 3537] = 0;
        memory[ 3538] = 0;
        memory[ 3539] = 0;
        memory[ 3540] = 0;
        memory[ 3541] = 0;
        memory[ 3542] = 0;
        memory[ 3543] = 0;
        memory[ 3544] = 0;
        memory[ 3545] = 0;
        memory[ 3546] = 0;
        memory[ 3547] = 0;
        memory[ 3548] = 1;
        memory[ 3549] = 0;
        memory[ 3550] = 0;
        memory[ 3551] = 0;
        memory[ 3552] = 0;
        memory[ 3553] = 0;
        memory[ 3554] = 0;
        memory[ 3555] = 0;
        memory[ 3556] = 0;
        memory[ 3557] = 0;
        memory[ 3558] = 0;
        memory[ 3559] = 0;
        memory[ 3560] = 0;
        memory[ 3561] = 0;
        memory[ 3562] = 0;
        memory[ 3563] = 0;
        memory[ 3564] = 0;
        memory[ 3565] = 0;
        memory[ 3566] = 0;
        memory[ 3567] = 0;
        memory[ 3568] = 0;
        memory[ 3569] = 0;
        memory[ 3570] = 0;
        memory[ 3571] = 0;
        memory[ 3572] = 0;
        memory[ 3573] = 1;
        memory[ 3574] = 0;
        memory[ 3575] = 0;
        memory[ 3576] = 0;
        memory[ 3577] = 0;
        memory[ 3578] = 0;
        memory[ 3579] = 0;
        memory[ 3580] = 0;
        memory[ 3581] = 1;
        memory[ 3582] = 0;
        memory[ 3583] = 0;
        memory[ 3584] = 0;
        memory[ 3585] = 0;
        memory[ 3586] = 0;
        memory[ 3587] = 0;
        memory[ 3588] = 0;
        memory[ 3589] = 0;
        memory[ 3590] = 0;
        memory[ 3591] = 0;
        memory[ 3592] = 0;
        memory[ 3593] = 1;
        memory[ 3594] = 0;
        memory[ 3595] = 0;
        memory[ 3596] = 0;
        memory[ 3597] = 0;
        memory[ 3598] = 0;
        memory[ 3599] = 0;
        memory[ 3600] = 0;
        memory[ 3601] = 0;
        memory[ 3602] = 0;
        memory[ 3603] = 0;
        memory[ 3604] = 0;
        memory[ 3605] = 0;
        memory[ 3606] = 0;
        memory[ 3607] = 0;
        memory[ 3608] = 0;
        memory[ 3609] = 0;
        memory[ 3610] = 1;
        memory[ 3611] = 0;
        memory[ 3612] = 0;
        memory[ 3613] = 0;
        memory[ 3614] = 0;
        memory[ 3615] = 0;
        memory[ 3616] = 0;
        memory[ 3617] = 0;
        memory[ 3618] = 0;
        memory[ 3619] = 0;
        memory[ 3620] = 0;
        memory[ 3621] = 0;
        memory[ 3622] = 0;
        memory[ 3623] = 0;
        memory[ 3624] = 0;
        memory[ 3625] = 0;
        memory[ 3626] = 0;
        memory[ 3627] = 0;
        memory[ 3628] = 0;
        memory[ 3629] = 0;
        memory[ 3630] = 0;
        memory[ 3631] = 0;
        memory[ 3632] = 0;
        memory[ 3633] = 0;
        memory[ 3634] = 0;
        memory[ 3635] = 1;
        memory[ 3636] = 0;
        memory[ 3637] = 0;
        memory[ 3638] = 0;
        memory[ 3639] = 0;
        memory[ 3640] = 0;
        memory[ 3641] = 0;
        memory[ 3642] = 0;
        memory[ 3643] = 0;
        memory[ 3644] = 0;
        memory[ 3645] = 0;
        memory[ 3646] = 0;
        memory[ 3647] = 0;
        memory[ 3648] = 0;
        memory[ 3649] = 0;
        memory[ 3650] = 0;
        memory[ 3651] = 0;
        memory[ 3652] = 0;
        memory[ 3653] = 0;
        memory[ 3654] = 0;
        memory[ 3655] = 0;
        memory[ 3656] = 0;
        memory[ 3657] = 0;
        memory[ 3658] = 0;
        memory[ 3659] = 0;
        memory[ 3660] = 0;
        memory[ 3661] = 0;
        memory[ 3662] = 0;
        memory[ 3663] = 0;
        memory[ 3664] = 0;
        memory[ 3665] = 0;
        memory[ 3666] = 0;
        memory[ 3667] = 1;
        memory[ 3668] = 0;
        memory[ 3669] = 0;
        memory[ 3670] = 0;
        memory[ 3671] = 0;
        memory[ 3672] = 0;
        memory[ 3673] = 0;
        memory[ 3674] = 0;
        memory[ 3675] = 0;
        memory[ 3676] = 0;
        memory[ 3677] = 0;
        memory[ 3678] = 1;
        memory[ 3679] = 0;
        memory[ 3680] = 0;
        memory[ 3681] = 0;
        memory[ 3682] = 0;
        memory[ 3683] = 0;
        memory[ 3684] = 0;
        memory[ 3685] = 0;
        memory[ 3686] = 0;
        memory[ 3687] = 0;
        memory[ 3688] = 0;
        memory[ 3689] = 1;
        memory[ 3690] = 0;
        memory[ 3691] = 0;
        memory[ 3692] = 0;
        memory[ 3693] = 1;
        memory[ 3694] = 1;
        memory[ 3695] = 0;
        memory[ 3696] = 0;
        memory[ 3697] = 0;
        memory[ 3698] = 0;
        memory[ 3699] = 1;
        memory[ 3700] = 0;
        memory[ 3701] = 0;
        memory[ 3702] = 0;
        memory[ 3703] = 0;
        memory[ 3704] = 0;
        memory[ 3705] = 0;
        memory[ 3706] = 1;
        memory[ 3707] = 0;
        memory[ 3708] = 0;
        memory[ 3709] = 0;
        memory[ 3710] = 0;
        memory[ 3711] = 0;
        memory[ 3712] = 0;
        memory[ 3713] = 0;
        memory[ 3714] = 0;
        memory[ 3715] = 0;
        memory[ 3716] = 0;
        memory[ 3717] = 0;
        memory[ 3718] = 0;
        memory[ 3719] = 0;
        memory[ 3720] = 0;
        memory[ 3721] = 0;
        memory[ 3722] = 0;
        memory[ 3723] = 0;
        memory[ 3724] = 0;
        memory[ 3725] = 1;
        memory[ 3726] = 1;
        memory[ 3727] = 0;
        memory[ 3728] = 0;
        memory[ 3729] = 0;
        memory[ 3730] = 0;
        memory[ 3731] = 0;
        memory[ 3732] = 0;
        memory[ 3733] = 0;
        memory[ 3734] = 0;
        memory[ 3735] = 0;
        memory[ 3736] = 0;
        memory[ 3737] = 0;
        memory[ 3738] = 0;
        memory[ 3739] = 0;
        memory[ 3740] = 0;
        memory[ 3741] = 0;
        memory[ 3742] = 0;
        memory[ 3743] = 0;
        memory[ 3744] = 0;
        memory[ 3745] = 0;
        memory[ 3746] = 0;
        memory[ 3747] = 0;
        memory[ 3748] = 0;
        memory[ 3749] = 0;
        memory[ 3750] = 0;
        memory[ 3751] = 0;
        memory[ 3752] = 0;
        memory[ 3753] = 0;
        memory[ 3754] = 0;
        memory[ 3755] = 0;
        memory[ 3756] = 0;
        memory[ 3757] = 0;
        memory[ 3758] = 0;
        memory[ 3759] = 0;
        memory[ 3760] = 0;
        memory[ 3761] = 0;
        memory[ 3762] = 0;
        memory[ 3763] = 0;
        memory[ 3764] = 0;
        memory[ 3765] = 1;
        memory[ 3766] = 1;
        memory[ 3767] = 1;
        memory[ 3768] = 0;
        memory[ 3769] = 0;
        memory[ 3770] = 0;
        memory[ 3771] = 0;
        memory[ 3772] = 0;
        memory[ 3773] = 0;
        memory[ 3774] = 0;
        memory[ 3775] = 0;
        memory[ 3776] = 0;
        memory[ 3777] = 0;
        memory[ 3778] = 0;
        memory[ 3779] = 0;
        memory[ 3780] = 0;
        memory[ 3781] = 1;
        memory[ 3782] = 0;
        memory[ 3783] = 1;
        memory[ 3784] = 1;
        memory[ 3785] = 0;
        memory[ 3786] = 0;
        memory[ 3787] = 0;
        memory[ 3788] = 0;
        memory[ 3789] = 0;
        memory[ 3790] = 0;
        memory[ 3791] = 0;
        memory[ 3792] = 0;
        memory[ 3793] = 0;
        memory[ 3794] = 1;
        memory[ 3795] = 0;
        memory[ 3796] = 0;
        memory[ 3797] = 0;
        memory[ 3798] = 0;
        memory[ 3799] = 0;
        memory[ 3800] = 0;
        memory[ 3801] = 0;
        memory[ 3802] = 0;
        memory[ 3803] = 0;
        memory[ 3804] = 0;
        memory[ 3805] = 0;
        memory[ 3806] = 0;
        memory[ 3807] = 0;
        memory[ 3808] = 0;
        memory[ 3809] = 0;
        memory[ 3810] = 0;
        memory[ 3811] = 0;
        memory[ 3812] = 1;
        memory[ 3813] = 1;
        memory[ 3814] = 1;
        memory[ 3815] = 0;
        memory[ 3816] = 0;
        memory[ 3817] = 0;
        memory[ 3818] = 0;
        memory[ 3819] = 0;
        memory[ 3820] = 0;
        memory[ 3821] = 0;
        memory[ 3822] = 0;
        memory[ 3823] = 0;
        memory[ 3824] = 0;
        memory[ 3825] = 0;
        memory[ 3826] = 0;
        memory[ 3827] = 0;
        memory[ 3828] = 0;
        memory[ 3829] = 0;
        memory[ 3830] = 0;
        memory[ 3831] = 0;
        memory[ 3832] = 0;
        memory[ 3833] = 1;
        memory[ 3834] = 1;
        memory[ 3835] = 0;
        memory[ 3836] = 0;
        memory[ 3837] = 0;
        memory[ 3838] = 0;
        memory[ 3839] = 0;
        memory[ 3840] = 0;
        memory[ 3841] = 0;
        memory[ 3842] = 0;
        memory[ 3843] = 0;
        memory[ 3844] = 0;
        memory[ 3845] = 0;
        memory[ 3846] = 0;
        memory[ 3847] = 0;
        memory[ 3848] = 0;
        memory[ 3849] = 0;
        memory[ 3850] = 0;
        memory[ 3851] = 0;
        memory[ 3852] = 0;
        memory[ 3853] = 0;
        memory[ 3854] = 0;
        memory[ 3855] = 1;
        memory[ 3856] = 0;
        memory[ 3857] = 0;
        memory[ 3858] = 0;
        memory[ 3859] = 0;
        memory[ 3860] = 0;
        memory[ 3861] = 0;
        memory[ 3862] = 0;
        memory[ 3863] = 0;
        memory[ 3864] = 0;
        memory[ 3865] = 0;
        memory[ 3866] = 0;
        memory[ 3867] = 0;
        memory[ 3868] = 1;
        memory[ 3869] = 0;
        memory[ 3870] = 0;
        memory[ 3871] = 1;
        memory[ 3872] = 0;
        memory[ 3873] = 0;
        memory[ 3874] = 0;
        memory[ 3875] = 0;
        memory[ 3876] = 0;
        memory[ 3877] = 0;
        memory[ 3878] = 0;
        memory[ 3879] = 0;
        memory[ 3880] = 0;
        memory[ 3881] = 0;
        memory[ 3882] = 0;
        memory[ 3883] = 0;
        memory[ 3884] = 0;
        memory[ 3885] = 0;
        memory[ 3886] = 0;
        memory[ 3887] = 0;
        memory[ 3888] = 0;
        memory[ 3889] = 0;
        memory[ 3890] = 0;
        memory[ 3891] = 0;
        memory[ 3892] = 0;
        memory[ 3893] = 1;
        memory[ 3894] = 1;
        memory[ 3895] = 1;
        memory[ 3896] = 1;
        memory[ 3897] = 1;
        memory[ 3898] = 0;
        memory[ 3899] = 0;
        memory[ 3900] = 0;
        memory[ 3901] = 0;
        memory[ 3902] = 0;
        memory[ 3903] = 0;
        memory[ 3904] = 0;
        memory[ 3905] = 0;
        memory[ 3906] = 0;
        memory[ 3907] = 0;
        memory[ 3908] = 0;
        memory[ 3909] = 0;
        memory[ 3910] = 0;
        memory[ 3911] = 0;
        memory[ 3912] = 0;
        memory[ 3913] = 0;
        memory[ 3914] = 0;
        memory[ 3915] = 0;
        memory[ 3916] = 0;
        memory[ 3917] = 1;
        memory[ 3918] = 1;
        memory[ 3919] = 1;
        memory[ 3920] = 0;
        memory[ 3921] = 0;
        memory[ 3922] = 0;
        memory[ 3923] = 0;
        memory[ 3924] = 0;
        memory[ 3925] = 0;
        memory[ 3926] = 0;
        memory[ 3927] = 0;
        memory[ 3928] = 0;
        memory[ 3929] = 0;
        memory[ 3930] = 0;
        memory[ 3931] = 0;
        memory[ 3932] = 0;
        memory[ 3933] = 0;
        memory[ 3934] = 0;
        memory[ 3935] = 1;
        memory[ 3936] = 1;
        memory[ 3937] = 0;
        memory[ 3938] = 0;
        memory[ 3939] = 0;
        memory[ 3940] = 0;
        memory[ 3941] = 0;
        memory[ 3942] = 0;
        memory[ 3943] = 0;
        memory[ 3944] = 1;
        memory[ 3945] = 1;
        memory[ 3946] = 1;
        memory[ 3947] = 0;
        memory[ 3948] = 0;
        memory[ 3949] = 1;
        memory[ 3950] = 1;
        memory[ 3951] = 1;
        memory[ 3952] = 0;
        memory[ 3953] = 0;
        memory[ 3954] = 0;
        memory[ 3955] = 0;
        memory[ 3956] = 0;
        memory[ 3957] = 0;
        memory[ 3958] = 0;
        memory[ 3959] = 1;
        memory[ 3960] = 1;
        memory[ 3961] = 0;
        memory[ 3962] = 0;
        memory[ 3963] = 0;
        memory[ 3964] = 0;
        memory[ 3965] = 0;
        memory[ 3966] = 0;
        memory[ 3967] = 0;
        memory[ 3968] = 0;
        memory[ 3969] = 0;
        memory[ 3970] = 0;
        memory[ 3971] = 0;
        memory[ 3972] = 0;
        memory[ 3973] = 0;
        memory[ 3974] = 0;
        memory[ 3975] = 0;
        memory[ 3976] = 0;
        memory[ 3977] = 0;
        memory[ 3978] = 0;
        memory[ 3979] = 0;
        memory[ 3980] = 0;
        memory[ 3981] = 1;
        memory[ 3982] = 0;
        memory[ 3983] = 0;
        memory[ 3984] = 0;
        memory[ 3985] = 0;
        memory[ 3986] = 0;
        memory[ 3987] = 0;
        memory[ 3988] = 0;
        memory[ 3989] = 0;
        memory[ 3990] = 0;
        memory[ 3991] = 0;
        memory[ 3992] = 0;
        memory[ 3993] = 0;
        memory[ 3994] = 0;
        memory[ 3995] = 0;
        memory[ 3996] = 0;
        memory[ 3997] = 0;
        memory[ 3998] = 0;
        memory[ 3999] = 0;
        memory[ 4000] = 0;
        memory[ 4001] = 1;
        memory[ 4002] = 0;
        memory[ 4003] = 0;
        memory[ 4004] = 0;
        memory[ 4005] = 0;
        memory[ 4006] = 0;
        memory[ 4007] = 0;
        memory[ 4008] = 1;
        memory[ 4009] = 0;
        memory[ 4010] = 0;
        memory[ 4011] = 0;
        memory[ 4012] = 0;
        memory[ 4013] = 0;
        memory[ 4014] = 0;
        memory[ 4015] = 0;
        memory[ 4016] = 0;
        memory[ 4017] = 0;
        memory[ 4018] = 0;
        memory[ 4019] = 1;
        memory[ 4020] = 1;
        memory[ 4021] = 0;
        memory[ 4022] = 0;
        memory[ 4023] = 0;
        memory[ 4024] = 0;
        memory[ 4025] = 0;
        memory[ 4026] = 0;
        memory[ 4027] = 0;
        memory[ 4028] = 0;
        memory[ 4029] = 0;
        memory[ 4030] = 0;
        memory[ 4031] = 0;
        memory[ 4032] = 0;
        memory[ 4033] = 0;
        memory[ 4034] = 0;
        memory[ 4035] = 0;
        memory[ 4036] = 0;
        memory[ 4037] = 1;
        memory[ 4038] = 0;
        memory[ 4039] = 0;
        memory[ 4040] = 0;
        memory[ 4041] = 0;
        memory[ 4042] = 0;
        memory[ 4043] = 0;
        memory[ 4044] = 0;
        memory[ 4045] = 1;
        memory[ 4046] = 0;
        memory[ 4047] = 0;
        memory[ 4048] = 1;
        memory[ 4049] = 0;
        memory[ 4050] = 0;
        memory[ 4051] = 0;
        memory[ 4052] = 0;
        memory[ 4053] = 0;
        memory[ 4054] = 0;
        memory[ 4055] = 0;
        memory[ 4056] = 0;
        memory[ 4057] = 0;
        memory[ 4058] = 0;
        memory[ 4059] = 0;
        memory[ 4060] = 0;
        memory[ 4061] = 0;
        memory[ 4062] = 1;
        memory[ 4063] = 1;
        memory[ 4064] = 1;
        memory[ 4065] = 0;
        memory[ 4066] = 1;
        memory[ 4067] = 1;
        memory[ 4068] = 0;
        memory[ 4069] = 0;
        memory[ 4070] = 0;
        memory[ 4071] = 0;
        memory[ 4072] = 0;
        memory[ 4073] = 0;
        memory[ 4074] = 0;
        memory[ 4075] = 0;
        memory[ 4076] = 0;
        memory[ 4077] = 0;
        memory[ 4078] = 0;
        memory[ 4079] = 0;
        memory[ 4080] = 0;
        memory[ 4081] = 0;
        memory[ 4082] = 0;
        memory[ 4083] = 0;
        memory[ 4084] = 0;
        memory[ 4085] = 0;
        memory[ 4086] = 0;
        memory[ 4087] = 0;
        memory[ 4088] = 0;
        memory[ 4089] = 0;
        memory[ 4090] = 0;
        memory[ 4091] = 0;
        memory[ 4092] = 0;
        memory[ 4093] = 0;
        memory[ 4094] = 0;
        memory[ 4095] = 0;
        memory[ 4096] = 1;
        memory[ 4097] = 0;
        memory[ 4098] = 1;
        memory[ 4099] = 1;
        memory[ 4100] = 0;
        memory[ 4101] = 0;
        memory[ 4102] = 1;
        memory[ 4103] = 0;
        memory[ 4104] = 0;
        memory[ 4105] = 0;
        memory[ 4106] = 0;
        memory[ 4107] = 1;
        memory[ 4108] = 1;
        memory[ 4109] = 0;
        memory[ 4110] = 0;
        memory[ 4111] = 0;
        memory[ 4112] = 0;
        memory[ 4113] = 0;
        memory[ 4114] = 0;
        memory[ 4115] = 0;
        memory[ 4116] = 0;
        memory[ 4117] = 0;
        memory[ 4118] = 0;
        memory[ 4119] = 0;
        memory[ 4120] = 0;
        memory[ 4121] = 0;
        memory[ 4122] = 0;
        memory[ 4123] = 0;
        memory[ 4124] = 0;
        memory[ 4125] = 0;
        memory[ 4126] = 0;
        memory[ 4127] = 0;
        memory[ 4128] = 0;
        memory[ 4129] = 0;
        memory[ 4130] = 0;
        memory[ 4131] = 0;
        memory[ 4132] = 0;
        memory[ 4133] = 0;
        memory[ 4134] = 1;
        memory[ 4135] = 0;
        memory[ 4136] = 0;
        memory[ 4137] = 1;
        memory[ 4138] = 0;
        memory[ 4139] = 0;
        memory[ 4140] = 0;
        memory[ 4141] = 1;
        memory[ 4142] = 1;
        memory[ 4143] = 0;
        memory[ 4144] = 0;
        memory[ 4145] = 1;
        memory[ 4146] = 0;
        memory[ 4147] = 0;
        memory[ 4148] = 0;
        memory[ 4149] = 0;
        memory[ 4150] = 1;
        memory[ 4151] = 1;
        memory[ 4152] = 0;
        memory[ 4153] = 0;
        memory[ 4154] = 1;
        memory[ 4155] = 0;
        memory[ 4156] = 0;
        memory[ 4157] = 0;
        memory[ 4158] = 0;
        memory[ 4159] = 0;
        memory[ 4160] = 0;
        memory[ 4161] = 0;
        memory[ 4162] = 0;
        memory[ 4163] = 0;
        memory[ 4164] = 0;
        memory[ 4165] = 0;
        memory[ 4166] = 0;
        memory[ 4167] = 0;
        memory[ 4168] = 0;
        memory[ 4169] = 0;
        memory[ 4170] = 0;
        memory[ 4171] = 0;
        memory[ 4172] = 0;
        memory[ 4173] = 0;
        memory[ 4174] = 0;
        memory[ 4175] = 0;
        memory[ 4176] = 0;
        memory[ 4177] = 0;
        memory[ 4178] = 0;
        memory[ 4179] = 0;
        memory[ 4180] = 0;
        memory[ 4181] = 0;
        memory[ 4182] = 0;
        memory[ 4183] = 0;
        memory[ 4184] = 0;
        memory[ 4185] = 0;
        memory[ 4186] = 0;
        memory[ 4187] = 0;
        memory[ 4188] = 0;
        memory[ 4189] = 0;
        memory[ 4190] = 1;
        memory[ 4191] = 1;
        memory[ 4192] = 0;
        memory[ 4193] = 0;
        memory[ 4194] = 0;
        memory[ 4195] = 1;
        memory[ 4196] = 0;
        memory[ 4197] = 1;
        memory[ 4198] = 1;
        memory[ 4199] = 0;
        memory[ 4200] = 0;
        memory[ 4201] = 0;
        memory[ 4202] = 0;
        memory[ 4203] = 0;
        memory[ 4204] = 0;
        memory[ 4205] = 0;
        memory[ 4206] = 0;
        memory[ 4207] = 0;
        memory[ 4208] = 0;
        memory[ 4209] = 0;
        memory[ 4210] = 0;
        memory[ 4211] = 0;
        memory[ 4212] = 0;
        memory[ 4213] = 0;
        memory[ 4214] = 0;
        memory[ 4215] = 0;
        memory[ 4216] = 0;
        memory[ 4217] = 1;
        memory[ 4218] = 0;
        memory[ 4219] = 0;
        memory[ 4220] = 0;
        memory[ 4221] = 0;
        memory[ 4222] = 0;
        memory[ 4223] = 0;
        memory[ 4224] = 0;
        memory[ 4225] = 0;
        memory[ 4226] = 0;
        memory[ 4227] = 1;
        memory[ 4228] = 0;
        memory[ 4229] = 0;
        memory[ 4230] = 0;
        memory[ 4231] = 0;
        memory[ 4232] = 0;
        memory[ 4233] = 0;
        memory[ 4234] = 0;
        memory[ 4235] = 0;
        memory[ 4236] = 1;
        memory[ 4237] = 0;
        memory[ 4238] = 0;
        memory[ 4239] = 0;
        memory[ 4240] = 0;
        memory[ 4241] = 0;
        memory[ 4242] = 0;
        memory[ 4243] = 0;
        memory[ 4244] = 0;
        memory[ 4245] = 0;
        memory[ 4246] = 0;
        memory[ 4247] = 0;
        memory[ 4248] = 0;
        memory[ 4249] = 0;
        memory[ 4250] = 0;
        memory[ 4251] = 0;
        memory[ 4252] = 0;
        memory[ 4253] = 0;
        memory[ 4254] = 0;
        memory[ 4255] = 0;
        memory[ 4256] = 0;
        memory[ 4257] = 0;
        memory[ 4258] = 0;
        memory[ 4259] = 0;
        memory[ 4260] = 0;
        memory[ 4261] = 0;
        memory[ 4262] = 0;
        memory[ 4263] = 0;
        memory[ 4264] = 0;
        memory[ 4265] = 0;
        memory[ 4266] = 0;
        memory[ 4267] = 0;
        memory[ 4268] = 0;
        memory[ 4269] = 0;
        memory[ 4270] = 0;
        memory[ 4271] = 0;
        memory[ 4272] = 0;
        memory[ 4273] = 1;
        memory[ 4274] = 0;
        memory[ 4275] = 0;
        memory[ 4276] = 0;
        memory[ 4277] = 0;
        memory[ 4278] = 0;
        memory[ 4279] = 0;
        memory[ 4280] = 0;
        memory[ 4281] = 1;
        memory[ 4282] = 1;
        memory[ 4283] = 1;
        memory[ 4284] = 0;
        memory[ 4285] = 0;
        memory[ 4286] = 0;
        memory[ 4287] = 0;
        memory[ 4288] = 0;
        memory[ 4289] = 0;
        memory[ 4290] = 0;
        memory[ 4291] = 0;
        memory[ 4292] = 1;
        memory[ 4293] = 1;
        memory[ 4294] = 0;
        memory[ 4295] = 0;
        memory[ 4296] = 0;
        memory[ 4297] = 1;
        memory[ 4298] = 1;
        memory[ 4299] = 0;
        memory[ 4300] = 0;
        memory[ 4301] = 0;
        memory[ 4302] = 1;
        memory[ 4303] = 0;
        memory[ 4304] = 0;
        memory[ 4305] = 0;
        memory[ 4306] = 0;
        memory[ 4307] = 0;
        memory[ 4308] = 0;
        memory[ 4309] = 0;
        memory[ 4310] = 0;
        memory[ 4311] = 0;
        memory[ 4312] = 1;
        memory[ 4313] = 1;
        memory[ 4314] = 0;
        memory[ 4315] = 0;
        memory[ 4316] = 1;
        memory[ 4317] = 0;
        memory[ 4318] = 0;
        memory[ 4319] = 0;
        memory[ 4320] = 0;
        memory[ 4321] = 0;
        memory[ 4322] = 0;
        memory[ 4323] = 0;
        memory[ 4324] = 0;
        memory[ 4325] = 1;
        memory[ 4326] = 0;
        memory[ 4327] = 0;
        memory[ 4328] = 1;
        memory[ 4329] = 1;
        memory[ 4330] = 1;
        memory[ 4331] = 0;
        memory[ 4332] = 0;
        memory[ 4333] = 0;
        memory[ 4334] = 0;
        memory[ 4335] = 0;
        memory[ 4336] = 0;
        memory[ 4337] = 1;
        memory[ 4338] = 0;
        memory[ 4339] = 0;
        memory[ 4340] = 0;
        memory[ 4341] = 0;
        memory[ 4342] = 0;
        memory[ 4343] = 0;
        memory[ 4344] = 0;
        memory[ 4345] = 0;
        memory[ 4346] = 0;
        memory[ 4347] = 0;
        memory[ 4348] = 0;
        memory[ 4349] = 0;
        memory[ 4350] = 0;
        memory[ 4351] = 0;
        memory[ 4352] = 0;
        memory[ 4353] = 0;
        memory[ 4354] = 0;
        memory[ 4355] = 0;
        memory[ 4356] = 0;
        memory[ 4357] = 0;
        memory[ 4358] = 0;
        memory[ 4359] = 0;
        memory[ 4360] = 0;
        memory[ 4361] = 0;
        memory[ 4362] = 1;
        memory[ 4363] = 0;
        memory[ 4364] = 0;
        memory[ 4365] = 0;
        memory[ 4366] = 0;
        memory[ 4367] = 0;
        memory[ 4368] = 0;
        memory[ 4369] = 0;
        memory[ 4370] = 1;
        memory[ 4371] = 0;
        memory[ 4372] = 0;
        memory[ 4373] = 0;
        memory[ 4374] = 0;
        memory[ 4375] = 1;
        memory[ 4376] = 1;
        memory[ 4377] = 0;
        memory[ 4378] = 0;
        memory[ 4379] = 0;
        memory[ 4380] = 0;
        memory[ 4381] = 0;
        memory[ 4382] = 0;
        memory[ 4383] = 0;
        memory[ 4384] = 0;
        memory[ 4385] = 1;
        memory[ 4386] = 1;
        memory[ 4387] = 1;
        memory[ 4388] = 0;
        memory[ 4389] = 0;
        memory[ 4390] = 0;
        memory[ 4391] = 0;
        memory[ 4392] = 0;
        memory[ 4393] = 0;
        memory[ 4394] = 0;
        memory[ 4395] = 0;
        memory[ 4396] = 0;
        memory[ 4397] = 0;
        memory[ 4398] = 1;
        memory[ 4399] = 0;
        memory[ 4400] = 0;
        memory[ 4401] = 0;
        memory[ 4402] = 0;
        memory[ 4403] = 1;
        memory[ 4404] = 0;
        memory[ 4405] = 0;
        memory[ 4406] = 0;
        memory[ 4407] = 0;
        memory[ 4408] = 0;
        memory[ 4409] = 0;
        memory[ 4410] = 0;
        memory[ 4411] = 0;
        memory[ 4412] = 0;
        memory[ 4413] = 0;
        memory[ 4414] = 0;
        memory[ 4415] = 0;
        memory[ 4416] = 0;
        memory[ 4417] = 0;
        memory[ 4418] = 0;
        memory[ 4419] = 0;
        memory[ 4420] = 0;
        memory[ 4421] = 0;
        memory[ 4422] = 0;
        memory[ 4423] = 0;
        memory[ 4424] = 0;
        memory[ 4425] = 0;
        memory[ 4426] = 1;
        memory[ 4427] = 1;
        memory[ 4428] = 1;
        memory[ 4429] = 0;
        memory[ 4430] = 0;
        memory[ 4431] = 0;
        memory[ 4432] = 0;
        memory[ 4433] = 0;
        memory[ 4434] = 0;
        memory[ 4435] = 0;
        memory[ 4436] = 0;
        memory[ 4437] = 0;
        memory[ 4438] = 0;
        memory[ 4439] = 0;
        memory[ 4440] = 0;
        memory[ 4441] = 0;
        memory[ 4442] = 1;
        memory[ 4443] = 0;
        memory[ 4444] = 0;
        memory[ 4445] = 0;
        memory[ 4446] = 0;
        memory[ 4447] = 0;
        memory[ 4448] = 0;
        memory[ 4449] = 0;
        memory[ 4450] = 0;
        memory[ 4451] = 0;
        memory[ 4452] = 1;
        memory[ 4453] = 0;
        memory[ 4454] = 0;
        memory[ 4455] = 0;
        memory[ 4456] = 0;
        memory[ 4457] = 1;
        memory[ 4458] = 0;
        memory[ 4459] = 1;
        memory[ 4460] = 1;
        memory[ 4461] = 0;
        memory[ 4462] = 0;
        memory[ 4463] = 0;
        memory[ 4464] = 0;
        memory[ 4465] = 0;
        memory[ 4466] = 1;
        memory[ 4467] = 0;
        memory[ 4468] = 0;
        memory[ 4469] = 0;
        memory[ 4470] = 0;
        memory[ 4471] = 0;
        memory[ 4472] = 0;
        memory[ 4473] = 0;
        memory[ 4474] = 0;
        memory[ 4475] = 1;
        memory[ 4476] = 0;
        memory[ 4477] = 0;
        memory[ 4478] = 0;
        memory[ 4479] = 0;
        memory[ 4480] = 0;
        memory[ 4481] = 0;
        memory[ 4482] = 0;
        memory[ 4483] = 0;
        memory[ 4484] = 0;
        memory[ 4485] = 1;
        memory[ 4486] = 0;
        memory[ 4487] = 0;
        memory[ 4488] = 0;
        memory[ 4489] = 0;
        memory[ 4490] = 0;
        memory[ 4491] = 0;
        memory[ 4492] = 0;
        memory[ 4493] = 0;
        memory[ 4494] = 0;
        memory[ 4495] = 0;
        memory[ 4496] = 0;
        memory[ 4497] = 0;
        memory[ 4498] = 0;
        memory[ 4499] = 0;
        memory[ 4500] = 0;
        memory[ 4501] = 1;
        memory[ 4502] = 1;
        memory[ 4503] = 0;
        memory[ 4504] = 0;
        memory[ 4505] = 1;
        memory[ 4506] = 0;
        memory[ 4507] = 0;
        memory[ 4508] = 0;
        memory[ 4509] = 0;
        memory[ 4510] = 0;
        memory[ 4511] = 0;
        memory[ 4512] = 1;
        memory[ 4513] = 0;
        memory[ 4514] = 0;
        memory[ 4515] = 0;
        memory[ 4516] = 0;
        memory[ 4517] = 0;
        memory[ 4518] = 0;
        memory[ 4519] = 0;
        memory[ 4520] = 0;
        memory[ 4521] = 0;
        memory[ 4522] = 0;
        memory[ 4523] = 0;
        memory[ 4524] = 0;
        memory[ 4525] = 1;
        memory[ 4526] = 0;
        memory[ 4527] = 0;
        memory[ 4528] = 0;
        memory[ 4529] = 0;
        memory[ 4530] = 1;
        memory[ 4531] = 1;
        memory[ 4532] = 0;
        memory[ 4533] = 0;
        memory[ 4534] = 0;
        memory[ 4535] = 0;
        memory[ 4536] = 0;
        memory[ 4537] = 0;
        memory[ 4538] = 0;
        memory[ 4539] = 0;
        memory[ 4540] = 0;
        memory[ 4541] = 0;
        memory[ 4542] = 0;
        memory[ 4543] = 0;
        memory[ 4544] = 0;
        memory[ 4545] = 0;
        memory[ 4546] = 0;
        memory[ 4547] = 0;
        memory[ 4548] = 0;
        memory[ 4549] = 0;
        memory[ 4550] = 0;
        memory[ 4551] = 0;
        memory[ 4552] = 0;
        memory[ 4553] = 0;
        memory[ 4554] = 0;
        memory[ 4555] = 0;
        memory[ 4556] = 0;
        memory[ 4557] = 0;
        memory[ 4558] = 0;
        memory[ 4559] = 0;
        memory[ 4560] = 0;
        memory[ 4561] = 0;
        memory[ 4562] = 0;
        memory[ 4563] = 0;
        memory[ 4564] = 0;
        memory[ 4565] = 1;
        memory[ 4566] = 0;
        memory[ 4567] = 0;
        memory[ 4568] = 0;
        memory[ 4569] = 0;
        memory[ 4570] = 0;
        memory[ 4571] = 1;
        memory[ 4572] = 0;
        memory[ 4573] = 0;
        memory[ 4574] = 0;
        memory[ 4575] = 0;
        memory[ 4576] = 0;
        memory[ 4577] = 0;
        memory[ 4578] = 0;
        memory[ 4579] = 0;
        memory[ 4580] = 0;
        memory[ 4581] = 0;
        memory[ 4582] = 1;
        memory[ 4583] = 1;
        memory[ 4584] = 0;
        memory[ 4585] = 0;
        memory[ 4586] = 0;
        memory[ 4587] = 0;
        memory[ 4588] = 0;
        memory[ 4589] = 0;
        memory[ 4590] = 0;
        memory[ 4591] = 0;
        memory[ 4592] = 0;
        memory[ 4593] = 0;
        memory[ 4594] = 0;
        memory[ 4595] = 0;
        memory[ 4596] = 0;
        memory[ 4597] = 0;
        memory[ 4598] = 0;
        memory[ 4599] = 0;
        memory[ 4600] = 0;
        memory[ 4601] = 0;
        memory[ 4602] = 1;
        memory[ 4603] = 0;
        memory[ 4604] = 0;
        memory[ 4605] = 0;
        memory[ 4606] = 1;
        memory[ 4607] = 0;
        memory[ 4608] = 0;
        memory[ 4609] = 0;
        memory[ 4610] = 1;
        memory[ 4611] = 1;
        memory[ 4612] = 1;
        memory[ 4613] = 1;
        memory[ 4614] = 1;
        memory[ 4615] = 0;
        memory[ 4616] = 0;
        memory[ 4617] = 0;
        memory[ 4618] = 0;
        memory[ 4619] = 0;
        memory[ 4620] = 0;
        memory[ 4621] = 0;
        memory[ 4622] = 0;
        memory[ 4623] = 1;
        memory[ 4624] = 0;
        memory[ 4625] = 0;
        memory[ 4626] = 0;
        memory[ 4627] = 0;
        memory[ 4628] = 0;
        memory[ 4629] = 0;
        memory[ 4630] = 0;
        memory[ 4631] = 0;
        memory[ 4632] = 1;
        memory[ 4633] = 0;
        memory[ 4634] = 0;
        memory[ 4635] = 0;
        memory[ 4636] = 0;
        memory[ 4637] = 0;
        memory[ 4638] = 0;
        memory[ 4639] = 0;
        memory[ 4640] = 0;
        memory[ 4641] = 0;
        memory[ 4642] = 0;
        memory[ 4643] = 0;
        memory[ 4644] = 0;
        memory[ 4645] = 0;
        memory[ 4646] = 1;
        memory[ 4647] = 0;
        memory[ 4648] = 0;
        memory[ 4649] = 0;
        memory[ 4650] = 0;
        memory[ 4651] = 0;
        memory[ 4652] = 0;
        memory[ 4653] = 0;
        memory[ 4654] = 1;
        memory[ 4655] = 0;
        memory[ 4656] = 0;
        memory[ 4657] = 0;
        memory[ 4658] = 0;
        memory[ 4659] = 0;
        memory[ 4660] = 0;
        memory[ 4661] = 0;
        memory[ 4662] = 0;
        memory[ 4663] = 0;
        memory[ 4664] = 0;
        memory[ 4665] = 0;
        memory[ 4666] = 0;
        memory[ 4667] = 0;
        memory[ 4668] = 1;
        memory[ 4669] = 0;
        memory[ 4670] = 0;
        memory[ 4671] = 0;
        memory[ 4672] = 0;
        memory[ 4673] = 0;
        memory[ 4674] = 0;
        memory[ 4675] = 0;
        memory[ 4676] = 0;
        memory[ 4677] = 0;
        memory[ 4678] = 0;
        memory[ 4679] = 1;
        memory[ 4680] = 0;
        memory[ 4681] = 0;
        memory[ 4682] = 0;
        memory[ 4683] = 0;
        memory[ 4684] = 0;
        memory[ 4685] = 0;
        memory[ 4686] = 0;
        memory[ 4687] = 0;
        memory[ 4688] = 1;
        memory[ 4689] = 0;
        memory[ 4690] = 0;
        memory[ 4691] = 1;
        memory[ 4692] = 1;
        memory[ 4693] = 0;
        memory[ 4694] = 0;
        memory[ 4695] = 1;
        memory[ 4696] = 1;
        memory[ 4697] = 0;
        memory[ 4698] = 0;
        memory[ 4699] = 0;
        memory[ 4700] = 1;
        memory[ 4701] = 0;
        memory[ 4702] = 0;
        memory[ 4703] = 0;
        memory[ 4704] = 0;
        memory[ 4705] = 0;
        memory[ 4706] = 0;
        memory[ 4707] = 0;
        memory[ 4708] = 1;
        memory[ 4709] = 0;
        memory[ 4710] = 0;
        memory[ 4711] = 0;
        memory[ 4712] = 0;
        memory[ 4713] = 0;
        memory[ 4714] = 0;
        memory[ 4715] = 0;
        memory[ 4716] = 0;
        memory[ 4717] = 0;
        memory[ 4718] = 0;
        memory[ 4719] = 0;
        memory[ 4720] = 0;
        memory[ 4721] = 0;
        memory[ 4722] = 0;
        memory[ 4723] = 0;
        memory[ 4724] = 0;
        memory[ 4725] = 0;
        memory[ 4726] = 0;
        memory[ 4727] = 1;
        memory[ 4728] = 1;
        memory[ 4729] = 0;
        memory[ 4730] = 0;
        memory[ 4731] = 0;
        memory[ 4732] = 0;
        memory[ 4733] = 1;
        memory[ 4734] = 1;
        memory[ 4735] = 0;
        memory[ 4736] = 0;
        memory[ 4737] = 0;
        memory[ 4738] = 0;
        memory[ 4739] = 0;
        memory[ 4740] = 0;
        memory[ 4741] = 0;
        memory[ 4742] = 0;
        memory[ 4743] = 0;
        memory[ 4744] = 0;
        memory[ 4745] = 0;
        memory[ 4746] = 0;
        memory[ 4747] = 0;
        memory[ 4748] = 1;
        memory[ 4749] = 0;
        memory[ 4750] = 0;
        memory[ 4751] = 0;
        memory[ 4752] = 0;
        memory[ 4753] = 0;
        memory[ 4754] = 0;
        memory[ 4755] = 0;
        memory[ 4756] = 0;
        memory[ 4757] = 0;
        memory[ 4758] = 0;
        memory[ 4759] = 1;
        memory[ 4760] = 1;
        memory[ 4761] = 0;
        memory[ 4762] = 0;
        memory[ 4763] = 0;
        memory[ 4764] = 0;
        memory[ 4765] = 0;
        memory[ 4766] = 0;
        memory[ 4767] = 0;
        memory[ 4768] = 0;
        memory[ 4769] = 0;
        memory[ 4770] = 0;
        memory[ 4771] = 0;
        memory[ 4772] = 0;
        memory[ 4773] = 0;
        memory[ 4774] = 0;
        memory[ 4775] = 0;
        memory[ 4776] = 0;
        memory[ 4777] = 0;
        memory[ 4778] = 0;
        memory[ 4779] = 0;
        memory[ 4780] = 1;
        memory[ 4781] = 1;
        memory[ 4782] = 1;
        memory[ 4783] = 1;
        memory[ 4784] = 0;
        memory[ 4785] = 0;
        memory[ 4786] = 0;
        memory[ 4787] = 0;
        memory[ 4788] = 0;
        memory[ 4789] = 0;
        memory[ 4790] = 0;
        memory[ 4791] = 0;
        memory[ 4792] = 0;
        memory[ 4793] = 0;
        memory[ 4794] = 0;
        memory[ 4795] = 0;
        memory[ 4796] = 0;
        memory[ 4797] = 0;
        memory[ 4798] = 0;
        memory[ 4799] = 0;
        memory[ 4800] = 0;
        memory[ 4801] = 0;
        memory[ 4802] = 0;
        memory[ 4803] = 0;
        memory[ 4804] = 0;
        memory[ 4805] = 0;
        memory[ 4806] = 0;
        memory[ 4807] = 0;
        memory[ 4808] = 0;
        memory[ 4809] = 0;
        memory[ 4810] = 0;
        memory[ 4811] = 0;
        memory[ 4812] = 0;
        memory[ 4813] = 0;
        memory[ 4814] = 0;
        memory[ 4815] = 0;
        memory[ 4816] = 0;
        memory[ 4817] = 0;
        memory[ 4818] = 0;
        memory[ 4819] = 0;
        memory[ 4820] = 0;
        memory[ 4821] = 0;
        memory[ 4822] = 0;
        memory[ 4823] = 0;
        memory[ 4824] = 0;
        memory[ 4825] = 0;
        memory[ 4826] = 0;
        memory[ 4827] = 0;
        memory[ 4828] = 0;
        memory[ 4829] = 0;
        memory[ 4830] = 0;
        memory[ 4831] = 0;
        memory[ 4832] = 0;
        memory[ 4833] = 1;
        memory[ 4834] = 1;
        memory[ 4835] = 0;
        memory[ 4836] = 0;
        memory[ 4837] = 0;
        memory[ 4838] = 0;
        memory[ 4839] = 0;
        memory[ 4840] = 0;
        memory[ 4841] = 0;
        memory[ 4842] = 0;
        memory[ 4843] = 0;
        memory[ 4844] = 0;
        memory[ 4845] = 1;
        memory[ 4846] = 0;
        memory[ 4847] = 0;
        memory[ 4848] = 0;
        memory[ 4849] = 0;
        memory[ 4850] = 0;
        memory[ 4851] = 0;
        memory[ 4852] = 0;
        memory[ 4853] = 0;
        memory[ 4854] = 0;
        memory[ 4855] = 1;
        memory[ 4856] = 1;
        memory[ 4857] = 1;
        memory[ 4858] = 0;
        memory[ 4859] = 0;
        memory[ 4860] = 0;
        memory[ 4861] = 1;
        memory[ 4862] = 0;
        memory[ 4863] = 0;
        memory[ 4864] = 0;
        memory[ 4865] = 0;
        memory[ 4866] = 0;
        memory[ 4867] = 0;
        memory[ 4868] = 0;
        memory[ 4869] = 0;
        memory[ 4870] = 0;
        memory[ 4871] = 1;
        memory[ 4872] = 0;
        memory[ 4873] = 0;
        memory[ 4874] = 0;
        memory[ 4875] = 0;
        memory[ 4876] = 0;
        memory[ 4877] = 0;
        memory[ 4878] = 0;
        memory[ 4879] = 0;
        memory[ 4880] = 0;
        memory[ 4881] = 0;
        memory[ 4882] = 0;
        memory[ 4883] = 0;
        memory[ 4884] = 0;
        memory[ 4885] = 0;
        memory[ 4886] = 0;
        memory[ 4887] = 0;
        memory[ 4888] = 0;
        memory[ 4889] = 0;
        memory[ 4890] = 0;
        memory[ 4891] = 0;
        memory[ 4892] = 0;
        memory[ 4893] = 0;
        memory[ 4894] = 0;
        memory[ 4895] = 0;
        memory[ 4896] = 0;
        memory[ 4897] = 0;
        memory[ 4898] = 0;
        memory[ 4899] = 0;
        memory[ 4900] = 0;
        memory[ 4901] = 0;
        memory[ 4902] = 0;
        memory[ 4903] = 0;
        memory[ 4904] = 1;
        memory[ 4905] = 1;
        memory[ 4906] = 0;
        memory[ 4907] = 0;
        memory[ 4908] = 0;
        memory[ 4909] = 0;
        memory[ 4910] = 0;
        memory[ 4911] = 0;
        memory[ 4912] = 0;
        memory[ 4913] = 0;
        memory[ 4914] = 0;
        memory[ 4915] = 0;
        memory[ 4916] = 0;
        memory[ 4917] = 0;
        memory[ 4918] = 0;
        memory[ 4919] = 0;
        memory[ 4920] = 0;
        memory[ 4921] = 0;
        memory[ 4922] = 0;
        memory[ 4923] = 0;
        memory[ 4924] = 0;
        memory[ 4925] = 1;
        memory[ 4926] = 0;
        memory[ 4927] = 0;
        memory[ 4928] = 0;
        memory[ 4929] = 0;
        memory[ 4930] = 0;
        memory[ 4931] = 0;
        memory[ 4932] = 0;
        memory[ 4933] = 0;
        memory[ 4934] = 0;
        memory[ 4935] = 1;
        memory[ 4936] = 1;
        memory[ 4937] = 0;
        memory[ 4938] = 0;
        memory[ 4939] = 0;
        memory[ 4940] = 0;
        memory[ 4941] = 0;
        memory[ 4942] = 0;
        memory[ 4943] = 1;
        memory[ 4944] = 1;
        memory[ 4945] = 0;
        memory[ 4946] = 0;
        memory[ 4947] = 0;
        memory[ 4948] = 0;
        memory[ 4949] = 0;
        memory[ 4950] = 0;
        memory[ 4951] = 0;
        memory[ 4952] = 0;
        memory[ 4953] = 0;
        memory[ 4954] = 1;
        memory[ 4955] = 0;
        memory[ 4956] = 0;
        memory[ 4957] = 0;
        memory[ 4958] = 1;
        memory[ 4959] = 1;
        memory[ 4960] = 0;
        memory[ 4961] = 0;
        memory[ 4962] = 0;
        memory[ 4963] = 0;
        memory[ 4964] = 1;
        memory[ 4965] = 0;
        memory[ 4966] = 1;
        memory[ 4967] = 0;
        memory[ 4968] = 0;
        memory[ 4969] = 0;
        memory[ 4970] = 0;
        memory[ 4971] = 0;
        memory[ 4972] = 0;
        memory[ 4973] = 0;
        memory[ 4974] = 0;
        memory[ 4975] = 0;
        memory[ 4976] = 0;
        memory[ 4977] = 0;
        memory[ 4978] = 0;
        memory[ 4979] = 0;
        memory[ 4980] = 0;
        memory[ 4981] = 0;
        memory[ 4982] = 0;
        memory[ 4983] = 0;
        memory[ 4984] = 0;
        memory[ 4985] = 0;
        memory[ 4986] = 0;
        memory[ 4987] = 0;
        memory[ 4988] = 0;
        memory[ 4989] = 0;
        memory[ 4990] = 0;
        memory[ 4991] = 0;
        memory[ 4992] = 0;
        memory[ 4993] = 1;
        memory[ 4994] = 0;
        memory[ 4995] = 0;
        memory[ 4996] = 0;
        memory[ 4997] = 0;
        memory[ 4998] = 0;
        memory[ 4999] = 0;
        memory[ 5000] = 0;
        memory[ 5001] = 0;
        memory[ 5002] = 0;
        memory[ 5003] = 0;
        memory[ 5004] = 0;
        memory[ 5005] = 0;
        memory[ 5006] = 0;
        memory[ 5007] = 0;
        memory[ 5008] = 0;
        memory[ 5009] = 0;
        memory[ 5010] = 0;
        memory[ 5011] = 0;
        memory[ 5012] = 0;
        memory[ 5013] = 0;
        memory[ 5014] = 0;
        memory[ 5015] = 0;
        memory[ 5016] = 0;
        memory[ 5017] = 0;
        memory[ 5018] = 0;
        memory[ 5019] = 0;
        memory[ 5020] = 0;
        memory[ 5021] = 0;
        memory[ 5022] = 0;
        memory[ 5023] = 0;
        memory[ 5024] = 0;
        memory[ 5025] = 0;
        memory[ 5026] = 0;
        memory[ 5027] = 0;
        memory[ 5028] = 0;
        memory[ 5029] = 0;
        memory[ 5030] = 1;
        memory[ 5031] = 0;
        memory[ 5032] = 0;
        memory[ 5033] = 0;
        memory[ 5034] = 0;
        memory[ 5035] = 0;
        memory[ 5036] = 0;
        memory[ 5037] = 0;
        memory[ 5038] = 0;
        memory[ 5039] = 0;
        memory[ 5040] = 0;
        memory[ 5041] = 0;
        memory[ 5042] = 0;
        memory[ 5043] = 0;
        memory[ 5044] = 0;
        memory[ 5045] = 0;
        memory[ 5046] = 0;
        memory[ 5047] = 1;
        memory[ 5048] = 0;
        memory[ 5049] = 0;
        memory[ 5050] = 0;
        memory[ 5051] = 0;
        memory[ 5052] = 0;
        memory[ 5053] = 0;
        memory[ 5054] = 0;
        memory[ 5055] = 0;
        memory[ 5056] = 0;
        memory[ 5057] = 0;
        memory[ 5058] = 0;
        memory[ 5059] = 0;
        memory[ 5060] = 0;
        memory[ 5061] = 0;
        memory[ 5062] = 0;
        memory[ 5063] = 0;
        memory[ 5064] = 0;
        memory[ 5065] = 0;
        memory[ 5066] = 0;
        memory[ 5067] = 0;
        memory[ 5068] = 1;
        memory[ 5069] = 0;
        memory[ 5070] = 0;
        memory[ 5071] = 0;
        memory[ 5072] = 0;
        memory[ 5073] = 0;
        memory[ 5074] = 0;
        memory[ 5075] = 1;
        memory[ 5076] = 0;
        memory[ 5077] = 0;
        memory[ 5078] = 0;
        memory[ 5079] = 0;
        memory[ 5080] = 0;
        memory[ 5081] = 0;
        memory[ 5082] = 0;
        memory[ 5083] = 0;
        memory[ 5084] = 0;
        memory[ 5085] = 0;
        memory[ 5086] = 0;
        memory[ 5087] = 0;
        memory[ 5088] = 0;
        memory[ 5089] = 0;
        memory[ 5090] = 0;
        memory[ 5091] = 0;
        memory[ 5092] = 0;
        memory[ 5093] = 0;
        memory[ 5094] = 1;
        memory[ 5095] = 0;
        memory[ 5096] = 0;
        memory[ 5097] = 0;
        memory[ 5098] = 0;
        memory[ 5099] = 0;
        memory[ 5100] = 0;
        memory[ 5101] = 0;
        memory[ 5102] = 0;
        memory[ 5103] = 0;
        memory[ 5104] = 0;
        memory[ 5105] = 0;
        memory[ 5106] = 0;
        memory[ 5107] = 0;
        memory[ 5108] = 0;
        memory[ 5109] = 0;
        memory[ 5110] = 0;
        memory[ 5111] = 0;
        memory[ 5112] = 0;
        memory[ 5113] = 1;
        memory[ 5114] = 1;
        memory[ 5115] = 1;
        memory[ 5116] = 1;
        memory[ 5117] = 1;
        memory[ 5118] = 0;
        memory[ 5119] = 0;
        memory[ 5120] = 0;
        memory[ 5121] = 0;
        memory[ 5122] = 0;
        memory[ 5123] = 0;
        memory[ 5124] = 0;
        memory[ 5125] = 1;
        memory[ 5126] = 0;
        memory[ 5127] = 0;
        memory[ 5128] = 1;
        memory[ 5129] = 0;
        memory[ 5130] = 0;
        memory[ 5131] = 0;
        memory[ 5132] = 0;
        memory[ 5133] = 0;
        memory[ 5134] = 0;
        memory[ 5135] = 0;
        memory[ 5136] = 0;
        memory[ 5137] = 0;
        memory[ 5138] = 0;
        memory[ 5139] = 0;
        memory[ 5140] = 0;
        memory[ 5141] = 0;
        memory[ 5142] = 0;
        memory[ 5143] = 0;
        memory[ 5144] = 0;
        memory[ 5145] = 0;
        memory[ 5146] = 0;
        memory[ 5147] = 0;
        memory[ 5148] = 0;
        memory[ 5149] = 0;
        memory[ 5150] = 1;
        memory[ 5151] = 0;
        memory[ 5152] = 0;
        memory[ 5153] = 0;
        memory[ 5154] = 0;
        memory[ 5155] = 0;
        memory[ 5156] = 0;
        memory[ 5157] = 0;
        memory[ 5158] = 0;
        memory[ 5159] = 0;
        memory[ 5160] = 0;
        memory[ 5161] = 0;
        memory[ 5162] = 0;
        memory[ 5163] = 0;
        memory[ 5164] = 0;
        memory[ 5165] = 0;
        memory[ 5166] = 0;
        memory[ 5167] = 0;
        memory[ 5168] = 0;
        memory[ 5169] = 0;
        memory[ 5170] = 0;
        memory[ 5171] = 1;
        memory[ 5172] = 0;
        memory[ 5173] = 0;
        memory[ 5174] = 0;
        memory[ 5175] = 0;
        memory[ 5176] = 0;
        memory[ 5177] = 0;
        memory[ 5178] = 0;
        memory[ 5179] = 0;
        memory[ 5180] = 1;
        memory[ 5181] = 1;
        memory[ 5182] = 0;
        memory[ 5183] = 0;
        memory[ 5184] = 0;
        memory[ 5185] = 0;
        memory[ 5186] = 0;
        memory[ 5187] = 1;
        memory[ 5188] = 0;
        memory[ 5189] = 0;
        memory[ 5190] = 0;
        memory[ 5191] = 0;
        memory[ 5192] = 0;
        memory[ 5193] = 0;
        memory[ 5194] = 0;
        memory[ 5195] = 0;
        memory[ 5196] = 0;
        memory[ 5197] = 0;
        memory[ 5198] = 0;
        memory[ 5199] = 0;
        memory[ 5200] = 0;
        memory[ 5201] = 0;
        memory[ 5202] = 0;
        memory[ 5203] = 0;
        memory[ 5204] = 0;
        memory[ 5205] = 0;
        memory[ 5206] = 0;
        memory[ 5207] = 0;
        memory[ 5208] = 0;
        memory[ 5209] = 0;
        memory[ 5210] = 0;
        memory[ 5211] = 0;
        memory[ 5212] = 0;
        memory[ 5213] = 0;
        memory[ 5214] = 0;
        memory[ 5215] = 0;
        memory[ 5216] = 0;
        memory[ 5217] = 0;
        memory[ 5218] = 1;
        memory[ 5219] = 1;
        memory[ 5220] = 0;
        memory[ 5221] = 0;
        memory[ 5222] = 0;
        memory[ 5223] = 0;
        memory[ 5224] = 0;
        memory[ 5225] = 0;
        memory[ 5226] = 0;
        memory[ 5227] = 0;
        memory[ 5228] = 0;
        memory[ 5229] = 0;
        memory[ 5230] = 0;
        memory[ 5231] = 0;
        memory[ 5232] = 1;
        memory[ 5233] = 0;
        memory[ 5234] = 0;
        memory[ 5235] = 0;
        memory[ 5236] = 0;
        memory[ 5237] = 0;
        memory[ 5238] = 0;
        memory[ 5239] = 0;
        memory[ 5240] = 0;
        memory[ 5241] = 0;
        memory[ 5242] = 0;
        memory[ 5243] = 0;
        memory[ 5244] = 0;
        memory[ 5245] = 0;
        memory[ 5246] = 0;
        memory[ 5247] = 0;
        memory[ 5248] = 1;
        memory[ 5249] = 0;
        memory[ 5250] = 0;
        memory[ 5251] = 0;
        memory[ 5252] = 0;
        memory[ 5253] = 0;
        memory[ 5254] = 0;
        memory[ 5255] = 0;
        memory[ 5256] = 0;
        memory[ 5257] = 0;
        memory[ 5258] = 1;
        memory[ 5259] = 0;
        memory[ 5260] = 0;
        memory[ 5261] = 0;
        memory[ 5262] = 0;
        memory[ 5263] = 0;
        memory[ 5264] = 0;
        memory[ 5265] = 0;
        memory[ 5266] = 0;
        memory[ 5267] = 0;
        memory[ 5268] = 0;
        memory[ 5269] = 0;
        memory[ 5270] = 0;
        memory[ 5271] = 0;
        memory[ 5272] = 0;
        memory[ 5273] = 0;
        memory[ 5274] = 0;
        memory[ 5275] = 0;
        memory[ 5276] = 0;
        memory[ 5277] = 0;
        memory[ 5278] = 0;
        memory[ 5279] = 0;
        memory[ 5280] = 0;
        memory[ 5281] = 0;
        memory[ 5282] = 0;
        memory[ 5283] = 0;
        memory[ 5284] = 0;
        memory[ 5285] = 0;
        memory[ 5286] = 0;
        memory[ 5287] = 1;
        memory[ 5288] = 0;
        memory[ 5289] = 0;
        memory[ 5290] = 0;
        memory[ 5291] = 0;
        memory[ 5292] = 0;
        memory[ 5293] = 0;
        memory[ 5294] = 0;
        memory[ 5295] = 0;
        memory[ 5296] = 0;
        memory[ 5297] = 1;
        memory[ 5298] = 0;
        memory[ 5299] = 0;
        memory[ 5300] = 0;
        memory[ 5301] = 0;
        memory[ 5302] = 0;
        memory[ 5303] = 0;
        memory[ 5304] = 1;
        memory[ 5305] = 1;
        memory[ 5306] = 0;
        memory[ 5307] = 0;
        memory[ 5308] = 0;
        memory[ 5309] = 0;
        memory[ 5310] = 0;
        memory[ 5311] = 0;
        memory[ 5312] = 0;
        memory[ 5313] = 0;
        memory[ 5314] = 0;
        memory[ 5315] = 0;
        memory[ 5316] = 0;
        memory[ 5317] = 0;
        memory[ 5318] = 0;
        memory[ 5319] = 0;
        memory[ 5320] = 0;
        memory[ 5321] = 0;
        memory[ 5322] = 0;
        memory[ 5323] = 0;
        memory[ 5324] = 0;
        memory[ 5325] = 0;
        memory[ 5326] = 0;
        memory[ 5327] = 0;
        memory[ 5328] = 1;
        memory[ 5329] = 0;
        memory[ 5330] = 0;
        memory[ 5331] = 0;
        memory[ 5332] = 0;
        memory[ 5333] = 0;
        memory[ 5334] = 0;
        memory[ 5335] = 1;
        memory[ 5336] = 0;
        memory[ 5337] = 0;
        memory[ 5338] = 0;
        memory[ 5339] = 0;
        memory[ 5340] = 0;
        memory[ 5341] = 0;
        memory[ 5342] = 0;
        memory[ 5343] = 0;
        memory[ 5344] = 0;
        memory[ 5345] = 0;
        memory[ 5346] = 0;
        memory[ 5347] = 0;
        memory[ 5348] = 0;
        memory[ 5349] = 0;
        memory[ 5350] = 0;
        memory[ 5351] = 0;
        memory[ 5352] = 0;
        memory[ 5353] = 0;
        memory[ 5354] = 0;
        memory[ 5355] = 0;
        memory[ 5356] = 0;
        memory[ 5357] = 0;
        memory[ 5358] = 0;
        memory[ 5359] = 0;
        memory[ 5360] = 0;
        memory[ 5361] = 0;
        memory[ 5362] = 1;
        memory[ 5363] = 0;
        memory[ 5364] = 0;
        memory[ 5365] = 0;
        memory[ 5366] = 0;
        memory[ 5367] = 0;
        memory[ 5368] = 0;
        memory[ 5369] = 0;
        memory[ 5370] = 0;
        memory[ 5371] = 0;
        memory[ 5372] = 0;
        memory[ 5373] = 0;
        memory[ 5374] = 0;
        memory[ 5375] = 0;
        memory[ 5376] = 0;
        memory[ 5377] = 0;
        memory[ 5378] = 0;
        memory[ 5379] = 0;
        memory[ 5380] = 0;
        memory[ 5381] = 0;
        memory[ 5382] = 0;
        memory[ 5383] = 0;
        memory[ 5384] = 0;
        memory[ 5385] = 0;
        memory[ 5386] = 0;
        memory[ 5387] = 0;
        memory[ 5388] = 0;
        memory[ 5389] = 0;
        memory[ 5390] = 0;
        memory[ 5391] = 1;
        memory[ 5392] = 1;
        memory[ 5393] = 0;
        memory[ 5394] = 0;
        memory[ 5395] = 0;
        memory[ 5396] = 0;
        memory[ 5397] = 0;
        memory[ 5398] = 0;
        memory[ 5399] = 0;
        memory[ 5400] = 1;
        memory[ 5401] = 0;
        memory[ 5402] = 0;
        memory[ 5403] = 0;
        memory[ 5404] = 0;
        memory[ 5405] = 0;
        memory[ 5406] = 0;
        memory[ 5407] = 0;
        memory[ 5408] = 0;
        memory[ 5409] = 0;
        memory[ 5410] = 0;
        memory[ 5411] = 0;
        memory[ 5412] = 0;
        memory[ 5413] = 0;
        memory[ 5414] = 0;
        memory[ 5415] = 0;
        memory[ 5416] = 0;
        memory[ 5417] = 0;
        memory[ 5418] = 0;
        memory[ 5419] = 0;
        memory[ 5420] = 0;
        memory[ 5421] = 0;
        memory[ 5422] = 0;
        memory[ 5423] = 0;
        memory[ 5424] = 0;
        memory[ 5425] = 1;
        memory[ 5426] = 0;
        memory[ 5427] = 0;
        memory[ 5428] = 0;
        memory[ 5429] = 0;
        memory[ 5430] = 0;
        memory[ 5431] = 0;
        memory[ 5432] = 0;
        memory[ 5433] = 0;
        memory[ 5434] = 0;
        memory[ 5435] = 0;
        memory[ 5436] = 0;
        memory[ 5437] = 0;
        memory[ 5438] = 0;
        memory[ 5439] = 0;
        memory[ 5440] = 0;
        memory[ 5441] = 0;
        memory[ 5442] = 0;
        memory[ 5443] = 0;
        memory[ 5444] = 1;
        memory[ 5445] = 0;
        memory[ 5446] = 0;
        memory[ 5447] = 0;
        memory[ 5448] = 0;
        memory[ 5449] = 0;
        memory[ 5450] = 1;
        memory[ 5451] = 0;
        memory[ 5452] = 0;
        memory[ 5453] = 0;
        memory[ 5454] = 0;
        memory[ 5455] = 0;
        memory[ 5456] = 0;
        memory[ 5457] = 0;
        memory[ 5458] = 0;
        memory[ 5459] = 0;
        memory[ 5460] = 0;
        memory[ 5461] = 0;
        memory[ 5462] = 0;
        memory[ 5463] = 0;
        memory[ 5464] = 0;
        memory[ 5465] = 0;
        memory[ 5466] = 0;
        memory[ 5467] = 0;
        memory[ 5468] = 0;
        memory[ 5469] = 0;
        memory[ 5470] = 0;
        memory[ 5471] = 0;
        memory[ 5472] = 0;
        memory[ 5473] = 0;
        memory[ 5474] = 0;
        memory[ 5475] = 0;
        memory[ 5476] = 0;
        memory[ 5477] = 0;
        memory[ 5478] = 0;
        memory[ 5479] = 0;
        memory[ 5480] = 0;
        memory[ 5481] = 0;
        memory[ 5482] = 0;
        memory[ 5483] = 0;
        memory[ 5484] = 1;
        memory[ 5485] = 1;
        memory[ 5486] = 0;
        memory[ 5487] = 0;
        memory[ 5488] = 0;
        memory[ 5489] = 0;
        memory[ 5490] = 0;
        memory[ 5491] = 0;
        memory[ 5492] = 0;
        memory[ 5493] = 0;
        memory[ 5494] = 0;
        memory[ 5495] = 0;
        memory[ 5496] = 0;
        memory[ 5497] = 0;
        memory[ 5498] = 0;
        memory[ 5499] = 0;
        memory[ 5500] = 0;
        memory[ 5501] = 0;
        memory[ 5502] = 0;
        memory[ 5503] = 0;
        memory[ 5504] = 0;
        memory[ 5505] = 0;
        memory[ 5506] = 0;
        memory[ 5507] = 0;
        memory[ 5508] = 0;
        memory[ 5509] = 0;
        memory[ 5510] = 0;
        memory[ 5511] = 0;
        memory[ 5512] = 0;
        memory[ 5513] = 0;
        memory[ 5514] = 0;
        memory[ 5515] = 0;
        memory[ 5516] = 0;
        memory[ 5517] = 0;
        memory[ 5518] = 0;
        memory[ 5519] = 0;
        memory[ 5520] = 0;
        memory[ 5521] = 0;
        memory[ 5522] = 0;
        memory[ 5523] = 0;
        memory[ 5524] = 0;
        memory[ 5525] = 0;
        memory[ 5526] = 0;
        memory[ 5527] = 0;
        memory[ 5528] = 0;
        memory[ 5529] = 0;
        memory[ 5530] = 0;
        memory[ 5531] = 0;
        memory[ 5532] = 0;
        memory[ 5533] = 0;
        memory[ 5534] = 0;
        memory[ 5535] = 0;
        memory[ 5536] = 0;
        memory[ 5537] = 1;
        memory[ 5538] = 0;
        memory[ 5539] = 0;
        memory[ 5540] = 1;
        memory[ 5541] = 0;
        memory[ 5542] = 0;
        memory[ 5543] = 0;
        memory[ 5544] = 0;
        memory[ 5545] = 0;
        memory[ 5546] = 0;
        memory[ 5547] = 0;
        memory[ 5548] = 0;
        memory[ 5549] = 0;
        memory[ 5550] = 0;
        memory[ 5551] = 0;
        memory[ 5552] = 0;
        memory[ 5553] = 0;
        memory[ 5554] = 0;
        memory[ 5555] = 0;
        memory[ 5556] = 0;
        memory[ 5557] = 1;
        memory[ 5558] = 0;
        memory[ 5559] = 0;
        memory[ 5560] = 0;
        memory[ 5561] = 0;
        memory[ 5562] = 0;
        memory[ 5563] = 0;
        memory[ 5564] = 0;
        memory[ 5565] = 0;
        memory[ 5566] = 0;
        memory[ 5567] = 0;
        memory[ 5568] = 0;
        memory[ 5569] = 0;
        memory[ 5570] = 0;
        memory[ 5571] = 0;
        memory[ 5572] = 0;
        memory[ 5573] = 1;
        memory[ 5574] = 0;
        memory[ 5575] = 0;
        memory[ 5576] = 1;
        memory[ 5577] = 0;
        memory[ 5578] = 0;
        memory[ 5579] = 0;
        memory[ 5580] = 1;
        memory[ 5581] = 0;
        memory[ 5582] = 0;
        memory[ 5583] = 0;
        memory[ 5584] = 0;
        memory[ 5585] = 0;
        memory[ 5586] = 0;
        memory[ 5587] = 0;
        memory[ 5588] = 0;
        memory[ 5589] = 0;
        memory[ 5590] = 0;
        memory[ 5591] = 0;
        memory[ 5592] = 0;
        memory[ 5593] = 0;
        memory[ 5594] = 0;
        memory[ 5595] = 0;
        memory[ 5596] = 0;
        memory[ 5597] = 0;
        memory[ 5598] = 0;
        memory[ 5599] = 0;
        memory[ 5600] = 0;
        memory[ 5601] = 0;
        memory[ 5602] = 0;
        memory[ 5603] = 1;
        memory[ 5604] = 0;
        memory[ 5605] = 0;
        memory[ 5606] = 0;
        memory[ 5607] = 0;
        memory[ 5608] = 0;
        memory[ 5609] = 0;
        memory[ 5610] = 0;
        memory[ 5611] = 0;
        memory[ 5612] = 0;
        memory[ 5613] = 0;
        memory[ 5614] = 0;
        memory[ 5615] = 0;
        memory[ 5616] = 0;
        memory[ 5617] = 0;
        memory[ 5618] = 0;
        memory[ 5619] = 0;
        memory[ 5620] = 0;
        memory[ 5621] = 0;
        memory[ 5622] = 0;
        memory[ 5623] = 0;
        memory[ 5624] = 0;
        memory[ 5625] = 0;
        memory[ 5626] = 0;
        memory[ 5627] = 0;
        memory[ 5628] = 0;
        memory[ 5629] = 0;
        memory[ 5630] = 0;
        memory[ 5631] = 0;
        memory[ 5632] = 0;
        memory[ 5633] = 0;
        memory[ 5634] = 0;
        memory[ 5635] = 0;
        memory[ 5636] = 0;
        memory[ 5637] = 1;
        memory[ 5638] = 0;
        memory[ 5639] = 0;
        memory[ 5640] = 0;
        memory[ 5641] = 0;
        memory[ 5642] = 0;
        memory[ 5643] = 0;
        memory[ 5644] = 0;
        memory[ 5645] = 0;
        memory[ 5646] = 0;
        memory[ 5647] = 0;
        memory[ 5648] = 0;
        memory[ 5649] = 0;
        memory[ 5650] = 0;
        memory[ 5651] = 0;
        memory[ 5652] = 0;
        memory[ 5653] = 0;
        memory[ 5654] = 0;
        memory[ 5655] = 0;
        memory[ 5656] = 0;
        memory[ 5657] = 0;
        memory[ 5658] = 0;
        memory[ 5659] = 0;
        memory[ 5660] = 0;
        memory[ 5661] = 0;
        memory[ 5662] = 0;
        memory[ 5663] = 0;
        memory[ 5664] = 0;
        memory[ 5665] = 0;
        memory[ 5666] = 0;
        memory[ 5667] = 0;
        memory[ 5668] = 0;
        memory[ 5669] = 0;
        memory[ 5670] = 0;
        memory[ 5671] = 0;
        memory[ 5672] = 0;
        memory[ 5673] = 0;
        memory[ 5674] = 0;
        memory[ 5675] = 0;
        memory[ 5676] = 0;
        memory[ 5677] = 0;
        memory[ 5678] = 0;
        memory[ 5679] = 0;
        memory[ 5680] = 0;
        memory[ 5681] = 0;
        memory[ 5682] = 0;
        memory[ 5683] = 0;
        memory[ 5684] = 0;
        memory[ 5685] = 1;
        memory[ 5686] = 0;
        memory[ 5687] = 0;
        memory[ 5688] = 0;
        memory[ 5689] = 0;
        memory[ 5690] = 0;
        memory[ 5691] = 0;
        memory[ 5692] = 0;
        memory[ 5693] = 0;
        memory[ 5694] = 0;
        memory[ 5695] = 0;
        memory[ 5696] = 0;
        memory[ 5697] = 0;
        memory[ 5698] = 0;
        memory[ 5699] = 0;
        memory[ 5700] = 0;
        memory[ 5701] = 0;
        memory[ 5702] = 0;
        memory[ 5703] = 0;
        memory[ 5704] = 0;
        memory[ 5705] = 0;
        memory[ 5706] = 0;
        memory[ 5707] = 0;
        memory[ 5708] = 0;
        memory[ 5709] = 0;
        memory[ 5710] = 1;
        memory[ 5711] = 0;
        memory[ 5712] = 0;
        memory[ 5713] = 0;
        memory[ 5714] = 0;
        memory[ 5715] = 0;
        memory[ 5716] = 0;
        memory[ 5717] = 0;
        memory[ 5718] = 1;
        memory[ 5719] = 0;
        memory[ 5720] = 0;
        memory[ 5721] = 0;
        memory[ 5722] = 0;
        memory[ 5723] = 0;
        memory[ 5724] = 0;
        memory[ 5725] = 0;
        memory[ 5726] = 0;
        memory[ 5727] = 0;
        memory[ 5728] = 1;
        memory[ 5729] = 1;
        memory[ 5730] = 0;
        memory[ 5731] = 0;
        memory[ 5732] = 0;
        memory[ 5733] = 0;
        memory[ 5734] = 0;
        memory[ 5735] = 0;
        memory[ 5736] = 0;
        memory[ 5737] = 0;
        memory[ 5738] = 1;
        memory[ 5739] = 1;
        memory[ 5740] = 1;
        memory[ 5741] = 0;
        memory[ 5742] = 0;
        memory[ 5743] = 0;
        memory[ 5744] = 0;
        memory[ 5745] = 0;
        memory[ 5746] = 0;
        memory[ 5747] = 0;
        memory[ 5748] = 1;
        memory[ 5749] = 0;
        memory[ 5750] = 0;
        memory[ 5751] = 0;
        memory[ 5752] = 0;
        memory[ 5753] = 0;
        memory[ 5754] = 0;
        memory[ 5755] = 1;
        memory[ 5756] = 1;
        memory[ 5757] = 0;
        memory[ 5758] = 0;
        memory[ 5759] = 0;
        memory[ 5760] = 0;
        memory[ 5761] = 0;
        memory[ 5762] = 0;
        memory[ 5763] = 0;
        memory[ 5764] = 0;
        memory[ 5765] = 0;
        memory[ 5766] = 0;
        memory[ 5767] = 0;
        memory[ 5768] = 0;
        memory[ 5769] = 0;
        memory[ 5770] = 0;
        memory[ 5771] = 0;
        memory[ 5772] = 0;
        memory[ 5773] = 0;
        memory[ 5774] = 0;
        memory[ 5775] = 0;
        memory[ 5776] = 0;
        memory[ 5777] = 0;
        memory[ 5778] = 0;
        memory[ 5779] = 0;
        memory[ 5780] = 0;
        memory[ 5781] = 1;
        memory[ 5782] = 0;
        memory[ 5783] = 0;
        memory[ 5784] = 0;
        memory[ 5785] = 0;
        memory[ 5786] = 0;
        memory[ 5787] = 1;
        memory[ 5788] = 0;
        memory[ 5789] = 0;
        memory[ 5790] = 1;
        memory[ 5791] = 0;
        memory[ 5792] = 0;
        memory[ 5793] = 0;
        memory[ 5794] = 0;
        memory[ 5795] = 0;
        memory[ 5796] = 0;
        memory[ 5797] = 0;
        memory[ 5798] = 0;
        memory[ 5799] = 0;
        memory[ 5800] = 0;
        memory[ 5801] = 0;
        memory[ 5802] = 0;
        memory[ 5803] = 0;
        memory[ 5804] = 0;
        memory[ 5805] = 0;
        memory[ 5806] = 1;
        memory[ 5807] = 0;
        memory[ 5808] = 0;
        memory[ 5809] = 0;
        memory[ 5810] = 0;
        memory[ 5811] = 0;
        memory[ 5812] = 0;
        memory[ 5813] = 0;
        memory[ 5814] = 0;
        memory[ 5815] = 0;
        memory[ 5816] = 0;
        memory[ 5817] = 0;
        memory[ 5818] = 0;
        memory[ 5819] = 0;
        memory[ 5820] = 0;
        memory[ 5821] = 0;
        memory[ 5822] = 0;
        memory[ 5823] = 0;
        memory[ 5824] = 0;
        memory[ 5825] = 0;
        memory[ 5826] = 0;
        memory[ 5827] = 0;
        memory[ 5828] = 0;
        memory[ 5829] = 0;
        memory[ 5830] = 0;
        memory[ 5831] = 0;
        memory[ 5832] = 1;
        memory[ 5833] = 1;
        memory[ 5834] = 0;
        memory[ 5835] = 0;
        memory[ 5836] = 0;
        memory[ 5837] = 0;
        memory[ 5838] = 0;
        memory[ 5839] = 0;
        memory[ 5840] = 0;
        memory[ 5841] = 1;
        memory[ 5842] = 0;
        memory[ 5843] = 0;
        memory[ 5844] = 0;
        memory[ 5845] = 0;
        memory[ 5846] = 0;
        memory[ 5847] = 0;
        memory[ 5848] = 0;
        memory[ 5849] = 0;
        memory[ 5850] = 0;
        memory[ 5851] = 0;
        memory[ 5852] = 0;
        memory[ 5853] = 0;
        memory[ 5854] = 0;
        memory[ 5855] = 0;
        memory[ 5856] = 0;
        memory[ 5857] = 0;
        memory[ 5858] = 1;
        memory[ 5859] = 0;
        memory[ 5860] = 0;
        memory[ 5861] = 0;
        memory[ 5862] = 0;
        memory[ 5863] = 0;
        memory[ 5864] = 0;
        memory[ 5865] = 0;
        memory[ 5866] = 0;
        memory[ 5867] = 0;
        memory[ 5868] = 0;
        memory[ 5869] = 1;
        memory[ 5870] = 0;
        memory[ 5871] = 0;
        memory[ 5872] = 0;
        memory[ 5873] = 0;
        memory[ 5874] = 0;
        memory[ 5875] = 0;
        memory[ 5876] = 0;
        memory[ 5877] = 0;
        memory[ 5878] = 0;
        memory[ 5879] = 0;
        memory[ 5880] = 0;
        memory[ 5881] = 0;
        memory[ 5882] = 0;
        memory[ 5883] = 0;
        memory[ 5884] = 0;
        memory[ 5885] = 0;
        memory[ 5886] = 0;
        memory[ 5887] = 0;
        memory[ 5888] = 0;
        memory[ 5889] = 0;
        memory[ 5890] = 0;
        memory[ 5891] = 0;
        memory[ 5892] = 1;
        memory[ 5893] = 0;
        memory[ 5894] = 0;
        memory[ 5895] = 0;
        memory[ 5896] = 0;
        memory[ 5897] = 0;
        memory[ 5898] = 0;
        memory[ 5899] = 0;
        memory[ 5900] = 0;
        memory[ 5901] = 0;
        memory[ 5902] = 0;
        memory[ 5903] = 0;
        memory[ 5904] = 0;
        memory[ 5905] = 0;
        memory[ 5906] = 0;
        memory[ 5907] = 0;
        memory[ 5908] = 1;
        memory[ 5909] = 1;
        memory[ 5910] = 1;
        memory[ 5911] = 0;
        memory[ 5912] = 0;
        memory[ 5913] = 0;
        memory[ 5914] = 0;
        memory[ 5915] = 1;
        memory[ 5916] = 1;
        memory[ 5917] = 0;
        memory[ 5918] = 0;
        memory[ 5919] = 0;
        memory[ 5920] = 0;
        memory[ 5921] = 0;
        memory[ 5922] = 0;
        memory[ 5923] = 0;
        memory[ 5924] = 0;
        memory[ 5925] = 0;
        memory[ 5926] = 0;
        memory[ 5927] = 1;
        memory[ 5928] = 0;
        memory[ 5929] = 0;
        memory[ 5930] = 0;
        memory[ 5931] = 0;
        memory[ 5932] = 0;
        memory[ 5933] = 0;
        memory[ 5934] = 0;
        memory[ 5935] = 0;
        memory[ 5936] = 0;
        memory[ 5937] = 0;
        memory[ 5938] = 0;
        memory[ 5939] = 0;
        memory[ 5940] = 0;
        memory[ 5941] = 0;
        memory[ 5942] = 0;
        memory[ 5943] = 0;
        memory[ 5944] = 0;
        memory[ 5945] = 0;
        memory[ 5946] = 0;
        memory[ 5947] = 0;
        memory[ 5948] = 1;
        memory[ 5949] = 0;
        memory[ 5950] = 0;
        memory[ 5951] = 0;
        memory[ 5952] = 0;
        memory[ 5953] = 0;
        memory[ 5954] = 0;
        memory[ 5955] = 0;
        memory[ 5956] = 0;
        memory[ 5957] = 0;
        memory[ 5958] = 0;
        memory[ 5959] = 0;
        memory[ 5960] = 0;
        memory[ 5961] = 0;
        memory[ 5962] = 0;
        memory[ 5963] = 0;
        memory[ 5964] = 0;
        memory[ 5965] = 0;
        memory[ 5966] = 0;
        memory[ 5967] = 0;
        memory[ 5968] = 0;
        memory[ 5969] = 0;
        memory[ 5970] = 0;
        memory[ 5971] = 0;
        memory[ 5972] = 0;
        memory[ 5973] = 0;
        memory[ 5974] = 0;
        memory[ 5975] = 0;
        memory[ 5976] = 0;
        memory[ 5977] = 0;
        memory[ 5978] = 0;
        memory[ 5979] = 0;
        memory[ 5980] = 0;
        memory[ 5981] = 0;
        memory[ 5982] = 0;
        memory[ 5983] = 0;
        memory[ 5984] = 0;
        memory[ 5985] = 0;
        memory[ 5986] = 0;
        memory[ 5987] = 0;
        memory[ 5988] = 0;
        memory[ 5989] = 0;
        memory[ 5990] = 0;
        memory[ 5991] = 0;
        memory[ 5992] = 0;
        memory[ 5993] = 0;
        memory[ 5994] = 0;
        memory[ 5995] = 0;
        memory[ 5996] = 0;
        memory[ 5997] = 0;
        memory[ 5998] = 0;
        memory[ 5999] = 0;
        memory[ 6000] = 1;
        memory[ 6001] = 0;
        memory[ 6002] = 0;
        memory[ 6003] = 0;
        memory[ 6004] = 0;
        memory[ 6005] = 0;
        memory[ 6006] = 0;
        memory[ 6007] = 0;
        memory[ 6008] = 0;
        memory[ 6009] = 0;
        memory[ 6010] = 0;
        memory[ 6011] = 0;
        memory[ 6012] = 0;
        memory[ 6013] = 0;
        memory[ 6014] = 0;
        memory[ 6015] = 0;
        memory[ 6016] = 0;
        memory[ 6017] = 0;
        memory[ 6018] = 1;
        memory[ 6019] = 0;
        memory[ 6020] = 0;
        memory[ 6021] = 0;
        memory[ 6022] = 0;
        memory[ 6023] = 0;
        memory[ 6024] = 0;
        memory[ 6025] = 0;
        memory[ 6026] = 0;
        memory[ 6027] = 0;
        memory[ 6028] = 0;
        memory[ 6029] = 0;
        memory[ 6030] = 0;
        memory[ 6031] = 0;
        memory[ 6032] = 0;
        memory[ 6033] = 0;
        memory[ 6034] = 0;
        memory[ 6035] = 0;
        memory[ 6036] = 0;
        memory[ 6037] = 0;
        memory[ 6038] = 0;
        memory[ 6039] = 0;
        memory[ 6040] = 0;
        memory[ 6041] = 0;
        memory[ 6042] = 0;
        memory[ 6043] = 0;
        memory[ 6044] = 0;
        memory[ 6045] = 0;
        memory[ 6046] = 0;
        memory[ 6047] = 0;
        memory[ 6048] = 0;
        memory[ 6049] = 0;
        memory[ 6050] = 0;
        memory[ 6051] = 0;
        memory[ 6052] = 0;
        memory[ 6053] = 0;
        memory[ 6054] = 0;
        memory[ 6055] = 0;
        memory[ 6056] = 0;
        memory[ 6057] = 0;
        memory[ 6058] = 0;
        memory[ 6059] = 0;
        memory[ 6060] = 0;
        memory[ 6061] = 0;
        memory[ 6062] = 0;
        memory[ 6063] = 0;
        memory[ 6064] = 0;
        memory[ 6065] = 0;
        memory[ 6066] = 1;
        memory[ 6067] = 1;
        memory[ 6068] = 0;
        memory[ 6069] = 0;
        memory[ 6070] = 0;
        memory[ 6071] = 0;
        memory[ 6072] = 0;
        memory[ 6073] = 0;
        memory[ 6074] = 0;
        memory[ 6075] = 0;
        memory[ 6076] = 0;
        memory[ 6077] = 0;
        memory[ 6078] = 0;
        memory[ 6079] = 0;
        memory[ 6080] = 0;
        memory[ 6081] = 0;
        memory[ 6082] = 0;
        memory[ 6083] = 0;
        memory[ 6084] = 0;
        memory[ 6085] = 0;
        memory[ 6086] = 0;
        memory[ 6087] = 0;
        memory[ 6088] = 0;
        memory[ 6089] = 0;
        memory[ 6090] = 1;
        memory[ 6091] = 0;
        memory[ 6092] = 0;
        memory[ 6093] = 0;
        memory[ 6094] = 0;
        memory[ 6095] = 0;
        memory[ 6096] = 0;
        memory[ 6097] = 0;
        memory[ 6098] = 0;
        memory[ 6099] = 0;
        memory[ 6100] = 0;
        memory[ 6101] = 0;
        memory[ 6102] = 1;
        memory[ 6103] = 0;
        memory[ 6104] = 0;
        memory[ 6105] = 0;
        memory[ 6106] = 0;
        memory[ 6107] = 0;
        memory[ 6108] = 0;
        memory[ 6109] = 0;
        memory[ 6110] = 0;
        memory[ 6111] = 0;
        memory[ 6112] = 0;
        memory[ 6113] = 0;
        memory[ 6114] = 1;
        memory[ 6115] = 0;
        memory[ 6116] = 0;
        memory[ 6117] = 1;
        memory[ 6118] = 1;
        memory[ 6119] = 0;
        memory[ 6120] = 0;
        memory[ 6121] = 0;
        memory[ 6122] = 0;
        memory[ 6123] = 0;
        memory[ 6124] = 0;
        memory[ 6125] = 0;
        memory[ 6126] = 0;
        memory[ 6127] = 0;
        memory[ 6128] = 0;
        memory[ 6129] = 0;
        memory[ 6130] = 0;
        memory[ 6131] = 1;
        memory[ 6132] = 0;
        memory[ 6133] = 0;
        memory[ 6134] = 1;
        memory[ 6135] = 0;
        memory[ 6136] = 0;
        memory[ 6137] = 0;
        memory[ 6138] = 0;
        memory[ 6139] = 0;
        memory[ 6140] = 0;
        memory[ 6141] = 0;
        memory[ 6142] = 0;
        memory[ 6143] = 0;
        memory[ 6144] = 0;
        memory[ 6145] = 0;
        memory[ 6146] = 0;
        memory[ 6147] = 0;
        memory[ 6148] = 0;
        memory[ 6149] = 0;
        memory[ 6150] = 0;
        memory[ 6151] = 0;
        memory[ 6152] = 0;
        memory[ 6153] = 0;
        memory[ 6154] = 0;
        memory[ 6155] = 0;
        memory[ 6156] = 0;
        memory[ 6157] = 0;
        memory[ 6158] = 0;
        memory[ 6159] = 0;
        memory[ 6160] = 0;
        memory[ 6161] = 0;
        memory[ 6162] = 0;
        memory[ 6163] = 0;
        memory[ 6164] = 0;
        memory[ 6165] = 1;
        memory[ 6166] = 1;
        memory[ 6167] = 0;
        memory[ 6168] = 0;
        memory[ 6169] = 0;
        memory[ 6170] = 0;
        memory[ 6171] = 0;
        memory[ 6172] = 0;
        memory[ 6173] = 0;
        memory[ 6174] = 0;
        memory[ 6175] = 0;
        memory[ 6176] = 0;
        memory[ 6177] = 0;
        memory[ 6178] = 0;
        memory[ 6179] = 0;
        memory[ 6180] = 0;
        memory[ 6181] = 0;
        memory[ 6182] = 0;
        memory[ 6183] = 0;
        memory[ 6184] = 0;
        memory[ 6185] = 0;
        memory[ 6186] = 0;
        memory[ 6187] = 0;
        memory[ 6188] = 0;
        memory[ 6189] = 0;
        memory[ 6190] = 0;
        memory[ 6191] = 0;
        memory[ 6192] = 0;
        memory[ 6193] = 0;
        memory[ 6194] = 0;
        memory[ 6195] = 0;
        memory[ 6196] = 0;
        memory[ 6197] = 0;
        memory[ 6198] = 0;
        memory[ 6199] = 0;
        memory[ 6200] = 0;
        memory[ 6201] = 0;
        memory[ 6202] = 0;
        memory[ 6203] = 0;
        memory[ 6204] = 0;
        memory[ 6205] = 0;
        memory[ 6206] = 0;
        memory[ 6207] = 0;
        memory[ 6208] = 0;
        memory[ 6209] = 0;
        memory[ 6210] = 1;
        memory[ 6211] = 0;
        memory[ 6212] = 0;
        memory[ 6213] = 0;
        memory[ 6214] = 1;
        memory[ 6215] = 0;
        memory[ 6216] = 0;
        memory[ 6217] = 0;
        memory[ 6218] = 0;
        memory[ 6219] = 0;
        memory[ 6220] = 0;
        memory[ 6221] = 0;
        memory[ 6222] = 0;
        memory[ 6223] = 0;
        memory[ 6224] = 0;
        memory[ 6225] = 0;
        memory[ 6226] = 0;
        memory[ 6227] = 1;
        memory[ 6228] = 0;
        memory[ 6229] = 0;
        memory[ 6230] = 0;
        memory[ 6231] = 0;
        memory[ 6232] = 0;
        memory[ 6233] = 0;
        memory[ 6234] = 0;
        memory[ 6235] = 0;
        memory[ 6236] = 0;
        memory[ 6237] = 0;
        memory[ 6238] = 0;
        memory[ 6239] = 0;
        memory[ 6240] = 0;
        memory[ 6241] = 0;
        memory[ 6242] = 0;
        memory[ 6243] = 0;
        memory[ 6244] = 0;
        memory[ 6245] = 0;
        memory[ 6246] = 0;
        memory[ 6247] = 0;
        memory[ 6248] = 0;
        memory[ 6249] = 0;
        memory[ 6250] = 1;
        memory[ 6251] = 0;
        memory[ 6252] = 0;
        memory[ 6253] = 0;
        memory[ 6254] = 1;
        memory[ 6255] = 0;
        memory[ 6256] = 0;
        memory[ 6257] = 1;
        memory[ 6258] = 1;
        memory[ 6259] = 1;
        memory[ 6260] = 0;
        memory[ 6261] = 0;
        memory[ 6262] = 0;
        memory[ 6263] = 0;
        memory[ 6264] = 0;
        memory[ 6265] = 0;
        memory[ 6266] = 0;
        memory[ 6267] = 0;
        memory[ 6268] = 0;
        memory[ 6269] = 0;
        memory[ 6270] = 0;
        memory[ 6271] = 0;
        memory[ 6272] = 1;
        memory[ 6273] = 0;
        memory[ 6274] = 0;
        memory[ 6275] = 0;
        memory[ 6276] = 0;
        memory[ 6277] = 0;
        memory[ 6278] = 1;
        memory[ 6279] = 0;
        memory[ 6280] = 0;
        memory[ 6281] = 0;
        memory[ 6282] = 0;
        memory[ 6283] = 0;
        memory[ 6284] = 0;
        memory[ 6285] = 0;
        memory[ 6286] = 1;
        memory[ 6287] = 0;
        memory[ 6288] = 0;
        memory[ 6289] = 0;
        memory[ 6290] = 0;
        memory[ 6291] = 0;
        memory[ 6292] = 0;
        memory[ 6293] = 0;
        memory[ 6294] = 0;
        memory[ 6295] = 0;
        memory[ 6296] = 0;
        memory[ 6297] = 1;
        memory[ 6298] = 0;
        memory[ 6299] = 0;
        memory[ 6300] = 1;
        memory[ 6301] = 0;
        memory[ 6302] = 0;
        memory[ 6303] = 0;
        memory[ 6304] = 0;
        memory[ 6305] = 0;
        memory[ 6306] = 0;
        memory[ 6307] = 0;
        memory[ 6308] = 0;
        memory[ 6309] = 0;
        memory[ 6310] = 0;
        memory[ 6311] = 1;
        memory[ 6312] = 0;
        memory[ 6313] = 0;
        memory[ 6314] = 0;
        memory[ 6315] = 0;
        memory[ 6316] = 0;
        memory[ 6317] = 1;
        memory[ 6318] = 0;
        memory[ 6319] = 0;
        memory[ 6320] = 0;
        memory[ 6321] = 0;
        memory[ 6322] = 0;
        memory[ 6323] = 0;
        memory[ 6324] = 0;
        memory[ 6325] = 0;
        memory[ 6326] = 0;
        memory[ 6327] = 0;
        memory[ 6328] = 0;
        memory[ 6329] = 0;
        memory[ 6330] = 0;
        memory[ 6331] = 0;
        memory[ 6332] = 0;
        memory[ 6333] = 0;
        memory[ 6334] = 1;
        memory[ 6335] = 0;
        memory[ 6336] = 0;
        memory[ 6337] = 0;
        memory[ 6338] = 1;
        memory[ 6339] = 0;
        memory[ 6340] = 0;
        memory[ 6341] = 0;
        memory[ 6342] = 0;
        memory[ 6343] = 0;
        memory[ 6344] = 0;
        memory[ 6345] = 0;
        memory[ 6346] = 0;
        memory[ 6347] = 0;
        memory[ 6348] = 0;
        memory[ 6349] = 0;
        memory[ 6350] = 0;
        memory[ 6351] = 1;
        memory[ 6352] = 1;
        memory[ 6353] = 0;
        memory[ 6354] = 0;
        memory[ 6355] = 0;
        memory[ 6356] = 0;
        memory[ 6357] = 0;
        memory[ 6358] = 0;
        memory[ 6359] = 0;
        memory[ 6360] = 0;
        memory[ 6361] = 0;
        memory[ 6362] = 0;
        memory[ 6363] = 1;
        memory[ 6364] = 0;
        memory[ 6365] = 0;
        memory[ 6366] = 0;
        memory[ 6367] = 0;
        memory[ 6368] = 0;
        memory[ 6369] = 0;
        memory[ 6370] = 0;
        memory[ 6371] = 0;
        memory[ 6372] = 0;
        memory[ 6373] = 0;
        memory[ 6374] = 1;
        memory[ 6375] = 1;
        memory[ 6376] = 0;
        memory[ 6377] = 0;
        memory[ 6378] = 0;
        memory[ 6379] = 1;
        memory[ 6380] = 0;
        memory[ 6381] = 0;
        memory[ 6382] = 1;
        memory[ 6383] = 1;
        memory[ 6384] = 0;
        memory[ 6385] = 0;
        memory[ 6386] = 0;
        memory[ 6387] = 0;
        memory[ 6388] = 0;
        memory[ 6389] = 0;
        memory[ 6390] = 0;
        memory[ 6391] = 1;
        memory[ 6392] = 1;
        memory[ 6393] = 0;
        memory[ 6394] = 0;
        memory[ 6395] = 1;
        memory[ 6396] = 1;
        memory[ 6397] = 0;
        memory[ 6398] = 0;
        memory[ 6399] = 0;
        memory[ 6400] = 1;
        memory[ 6401] = 0;
        memory[ 6402] = 0;
        memory[ 6403] = 1;
        memory[ 6404] = 0;
        memory[ 6405] = 0;
        memory[ 6406] = 0;
        memory[ 6407] = 0;
        memory[ 6408] = 0;
        memory[ 6409] = 0;
        memory[ 6410] = 1;
        memory[ 6411] = 0;
        memory[ 6412] = 1;
        memory[ 6413] = 0;
        memory[ 6414] = 0;
        memory[ 6415] = 1;
        memory[ 6416] = 0;
        memory[ 6417] = 1;
        memory[ 6418] = 0;
        memory[ 6419] = 0;
        memory[ 6420] = 0;
        memory[ 6421] = 0;
        memory[ 6422] = 1;
        memory[ 6423] = 0;
        memory[ 6424] = 0;
        memory[ 6425] = 1;
        memory[ 6426] = 1;
        memory[ 6427] = 1;
        memory[ 6428] = 0;
        memory[ 6429] = 0;
        memory[ 6430] = 0;
        memory[ 6431] = 1;
        memory[ 6432] = 0;
        memory[ 6433] = 0;
        memory[ 6434] = 0;
        memory[ 6435] = 0;
        memory[ 6436] = 0;
        memory[ 6437] = 0;
        memory[ 6438] = 0;
        memory[ 6439] = 0;
        memory[ 6440] = 0;
        memory[ 6441] = 0;
        memory[ 6442] = 0;
        memory[ 6443] = 0;
        memory[ 6444] = 1;
        memory[ 6445] = 1;
        memory[ 6446] = 0;
        memory[ 6447] = 0;
        memory[ 6448] = 0;
        memory[ 6449] = 0;
        memory[ 6450] = 0;
        memory[ 6451] = 0;
        memory[ 6452] = 0;
        memory[ 6453] = 0;
        memory[ 6454] = 1;
        memory[ 6455] = 1;
        memory[ 6456] = 1;
        memory[ 6457] = 0;
        memory[ 6458] = 0;
        memory[ 6459] = 0;
        memory[ 6460] = 0;
        memory[ 6461] = 0;
        memory[ 6462] = 0;
        memory[ 6463] = 0;
        memory[ 6464] = 0;
        memory[ 6465] = 0;
        memory[ 6466] = 0;
        memory[ 6467] = 0;
        memory[ 6468] = 0;
        memory[ 6469] = 0;
        memory[ 6470] = 0;
        memory[ 6471] = 0;
        memory[ 6472] = 0;
        memory[ 6473] = 0;
        memory[ 6474] = 0;
        memory[ 6475] = 0;
        memory[ 6476] = 0;
        memory[ 6477] = 0;
        memory[ 6478] = 0;
        memory[ 6479] = 0;
        memory[ 6480] = 0;
        memory[ 6481] = 0;
        memory[ 6482] = 0;
        memory[ 6483] = 1;
        memory[ 6484] = 1;
        memory[ 6485] = 1;
        memory[ 6486] = 0;
        memory[ 6487] = 0;
        memory[ 6488] = 0;
        memory[ 6489] = 0;
        memory[ 6490] = 0;
        memory[ 6491] = 0;
        memory[ 6492] = 0;
        memory[ 6493] = 0;
        memory[ 6494] = 0;
        memory[ 6495] = 0;
        memory[ 6496] = 0;
        memory[ 6497] = 0;
        memory[ 6498] = 0;
        memory[ 6499] = 0;
        memory[ 6500] = 0;
        memory[ 6501] = 0;
        memory[ 6502] = 0;
        memory[ 6503] = 0;
        memory[ 6504] = 0;
        memory[ 6505] = 0;
        memory[ 6506] = 0;
        memory[ 6507] = 0;
        memory[ 6508] = 0;
        memory[ 6509] = 0;
        memory[ 6510] = 1;
        memory[ 6511] = 1;
        memory[ 6512] = 0;
        memory[ 6513] = 1;
        memory[ 6514] = 0;
        memory[ 6515] = 0;
        memory[ 6516] = 0;
        memory[ 6517] = 0;
        memory[ 6518] = 0;
        memory[ 6519] = 1;
        memory[ 6520] = 0;
        memory[ 6521] = 0;
        memory[ 6522] = 1;
        memory[ 6523] = 0;
        memory[ 6524] = 0;
        memory[ 6525] = 0;
        memory[ 6526] = 0;
        memory[ 6527] = 0;
        memory[ 6528] = 1;
        memory[ 6529] = 1;
        memory[ 6530] = 0;
        memory[ 6531] = 0;
        memory[ 6532] = 0;
        memory[ 6533] = 1;
        memory[ 6534] = 0;
        memory[ 6535] = 0;
        memory[ 6536] = 0;
        memory[ 6537] = 0;
        memory[ 6538] = 0;
        memory[ 6539] = 0;
        memory[ 6540] = 0;
        memory[ 6541] = 1;
        memory[ 6542] = 0;
        memory[ 6543] = 0;
        memory[ 6544] = 0;
        memory[ 6545] = 0;
        memory[ 6546] = 1;
        memory[ 6547] = 0;
        memory[ 6548] = 0;
        memory[ 6549] = 0;
        memory[ 6550] = 0;
        memory[ 6551] = 0;
        memory[ 6552] = 0;
        memory[ 6553] = 0;
        memory[ 6554] = 0;
        memory[ 6555] = 0;
        memory[ 6556] = 0;
        memory[ 6557] = 0;
        memory[ 6558] = 0;
        memory[ 6559] = 1;
        memory[ 6560] = 0;
        memory[ 6561] = 0;
        memory[ 6562] = 1;
        memory[ 6563] = 0;
        memory[ 6564] = 0;
        memory[ 6565] = 0;
        memory[ 6566] = 0;
        memory[ 6567] = 1;
        memory[ 6568] = 0;
        memory[ 6569] = 0;
        memory[ 6570] = 0;
        memory[ 6571] = 0;
        memory[ 6572] = 0;
        memory[ 6573] = 0;
        memory[ 6574] = 0;
        memory[ 6575] = 0;
        memory[ 6576] = 0;
        memory[ 6577] = 0;
        memory[ 6578] = 0;
        memory[ 6579] = 0;
        memory[ 6580] = 0;
        memory[ 6581] = 0;
        memory[ 6582] = 0;
        memory[ 6583] = 0;
        memory[ 6584] = 0;
        memory[ 6585] = 0;
        memory[ 6586] = 0;
        memory[ 6587] = 0;
        memory[ 6588] = 0;
        memory[ 6589] = 0;
        memory[ 6590] = 0;
        memory[ 6591] = 0;
        memory[ 6592] = 0;
        memory[ 6593] = 0;
        memory[ 6594] = 0;
        memory[ 6595] = 0;
        memory[ 6596] = 1;
        memory[ 6597] = 0;
        memory[ 6598] = 0;
        memory[ 6599] = 0;
        memory[ 6600] = 1;
        memory[ 6601] = 0;
        memory[ 6602] = 0;
        memory[ 6603] = 0;
        memory[ 6604] = 0;
        memory[ 6605] = 0;
        memory[ 6606] = 0;
        memory[ 6607] = 1;
        memory[ 6608] = 0;
        memory[ 6609] = 0;
        memory[ 6610] = 0;
        memory[ 6611] = 0;
        memory[ 6612] = 0;
        memory[ 6613] = 0;
        memory[ 6614] = 0;
        memory[ 6615] = 0;
        memory[ 6616] = 1;
        memory[ 6617] = 1;
        memory[ 6618] = 0;
        memory[ 6619] = 0;
        memory[ 6620] = 0;
        memory[ 6621] = 0;
        memory[ 6622] = 0;
        memory[ 6623] = 0;
        memory[ 6624] = 0;
        memory[ 6625] = 0;
        memory[ 6626] = 0;
        memory[ 6627] = 0;
        memory[ 6628] = 0;
        memory[ 6629] = 0;
        memory[ 6630] = 0;
        memory[ 6631] = 0;
        memory[ 6632] = 0;
        memory[ 6633] = 0;
        memory[ 6634] = 0;
        memory[ 6635] = 0;
        memory[ 6636] = 0;
        memory[ 6637] = 0;
        memory[ 6638] = 0;
        memory[ 6639] = 0;
        memory[ 6640] = 0;
        memory[ 6641] = 0;
        memory[ 6642] = 0;
        memory[ 6643] = 0;
        memory[ 6644] = 1;
        memory[ 6645] = 1;
        memory[ 6646] = 1;
        memory[ 6647] = 1;
        memory[ 6648] = 0;
        memory[ 6649] = 0;
        memory[ 6650] = 0;
        memory[ 6651] = 0;
        memory[ 6652] = 0;
        memory[ 6653] = 0;
        memory[ 6654] = 0;
        memory[ 6655] = 0;
        memory[ 6656] = 0;
        memory[ 6657] = 0;
        memory[ 6658] = 0;
        memory[ 6659] = 0;
        memory[ 6660] = 0;
        memory[ 6661] = 0;
        memory[ 6662] = 0;
        memory[ 6663] = 0;
        memory[ 6664] = 0;
        memory[ 6665] = 0;
        memory[ 6666] = 0;
        memory[ 6667] = 0;
        memory[ 6668] = 0;
        memory[ 6669] = 0;
        memory[ 6670] = 0;
        memory[ 6671] = 1;
        memory[ 6672] = 0;
        memory[ 6673] = 0;
        memory[ 6674] = 0;
        memory[ 6675] = 0;
        memory[ 6676] = 1;
        memory[ 6677] = 0;
        memory[ 6678] = 0;
        memory[ 6679] = 0;
        memory[ 6680] = 0;
        memory[ 6681] = 0;
        memory[ 6682] = 0;
        memory[ 6683] = 0;
        memory[ 6684] = 0;
        memory[ 6685] = 0;
        memory[ 6686] = 0;
        memory[ 6687] = 0;
        memory[ 6688] = 0;
        memory[ 6689] = 0;
        memory[ 6690] = 0;
        memory[ 6691] = 0;
        memory[ 6692] = 0;
        memory[ 6693] = 1;
        memory[ 6694] = 0;
        memory[ 6695] = 0;
        memory[ 6696] = 0;
        memory[ 6697] = 0;
        memory[ 6698] = 1;
        memory[ 6699] = 0;
        memory[ 6700] = 0;
        memory[ 6701] = 1;
        memory[ 6702] = 0;
        memory[ 6703] = 0;
        memory[ 6704] = 0;
        memory[ 6705] = 0;
        memory[ 6706] = 1;
        memory[ 6707] = 0;
        memory[ 6708] = 1;
        memory[ 6709] = 0;
        memory[ 6710] = 0;
        memory[ 6711] = 1;
        memory[ 6712] = 0;
        memory[ 6713] = 0;
        memory[ 6714] = 0;
        memory[ 6715] = 0;
        memory[ 6716] = 0;
        memory[ 6717] = 1;
        memory[ 6718] = 0;
        memory[ 6719] = 0;
        memory[ 6720] = 0;
        memory[ 6721] = 0;
        memory[ 6722] = 0;
        memory[ 6723] = 0;
        memory[ 6724] = 0;
        memory[ 6725] = 0;
        memory[ 6726] = 0;
        memory[ 6727] = 0;
        memory[ 6728] = 1;
        memory[ 6729] = 0;
        memory[ 6730] = 0;
        memory[ 6731] = 0;
        memory[ 6732] = 0;
        memory[ 6733] = 0;
        memory[ 6734] = 1;
        memory[ 6735] = 0;
        memory[ 6736] = 0;
        memory[ 6737] = 0;
        memory[ 6738] = 0;
        memory[ 6739] = 0;
        memory[ 6740] = 0;
        memory[ 6741] = 0;
        memory[ 6742] = 0;
        memory[ 6743] = 0;
        memory[ 6744] = 0;
        memory[ 6745] = 0;
        memory[ 6746] = 0;
        memory[ 6747] = 0;
        memory[ 6748] = 0;
        memory[ 6749] = 0;
        memory[ 6750] = 0;
        memory[ 6751] = 0;
        memory[ 6752] = 0;
        memory[ 6753] = 0;
        memory[ 6754] = 0;
        memory[ 6755] = 0;
        memory[ 6756] = 1;
        memory[ 6757] = 0;
        memory[ 6758] = 1;
        memory[ 6759] = 0;
        memory[ 6760] = 0;
        memory[ 6761] = 0;
        memory[ 6762] = 0;
        memory[ 6763] = 0;
        memory[ 6764] = 0;
        memory[ 6765] = 0;
        memory[ 6766] = 0;
        memory[ 6767] = 0;
        memory[ 6768] = 1;
        memory[ 6769] = 0;
        memory[ 6770] = 0;
        memory[ 6771] = 0;
        memory[ 6772] = 0;
        memory[ 6773] = 0;
        memory[ 6774] = 0;
        memory[ 6775] = 0;
        memory[ 6776] = 0;
        memory[ 6777] = 0;
        memory[ 6778] = 0;
        memory[ 6779] = 0;
        memory[ 6780] = 0;
        memory[ 6781] = 0;
        memory[ 6782] = 0;
        memory[ 6783] = 0;
        memory[ 6784] = 0;
        memory[ 6785] = 0;
        memory[ 6786] = 1;
        memory[ 6787] = 0;
        memory[ 6788] = 0;
        memory[ 6789] = 1;
        memory[ 6790] = 0;
        memory[ 6791] = 0;
        memory[ 6792] = 0;
        memory[ 6793] = 0;
        memory[ 6794] = 0;
        memory[ 6795] = 0;
        memory[ 6796] = 1;
        memory[ 6797] = 0;
        memory[ 6798] = 0;
        memory[ 6799] = 0;
        memory[ 6800] = 0;
        memory[ 6801] = 0;
        memory[ 6802] = 0;
        memory[ 6803] = 0;
        memory[ 6804] = 0;
        memory[ 6805] = 1;
        memory[ 6806] = 1;
        memory[ 6807] = 0;
        memory[ 6808] = 0;
        memory[ 6809] = 0;
        memory[ 6810] = 0;
        memory[ 6811] = 0;
        memory[ 6812] = 1;
        memory[ 6813] = 0;
        memory[ 6814] = 1;
        memory[ 6815] = 0;
        memory[ 6816] = 0;
        memory[ 6817] = 0;
        memory[ 6818] = 1;
        memory[ 6819] = 0;
        memory[ 6820] = 0;
        memory[ 6821] = 1;
        memory[ 6822] = 1;
        memory[ 6823] = 1;
        memory[ 6824] = 1;
        memory[ 6825] = 0;
        memory[ 6826] = 0;
        memory[ 6827] = 0;
        memory[ 6828] = 0;
        memory[ 6829] = 0;
        memory[ 6830] = 0;
        memory[ 6831] = 0;
        memory[ 6832] = 0;
        memory[ 6833] = 0;
        memory[ 6834] = 0;
        memory[ 6835] = 0;
        memory[ 6836] = 0;
        memory[ 6837] = 0;
        memory[ 6838] = 0;
        memory[ 6839] = 0;
        memory[ 6840] = 0;
        memory[ 6841] = 0;
        memory[ 6842] = 0;
        memory[ 6843] = 0;
        memory[ 6844] = 0;
        memory[ 6845] = 0;
        memory[ 6846] = 0;
        memory[ 6847] = 0;
        memory[ 6848] = 0;
        memory[ 6849] = 0;
        memory[ 6850] = 0;
        memory[ 6851] = 0;
        memory[ 6852] = 0;
        memory[ 6853] = 1;
        memory[ 6854] = 0;
        memory[ 6855] = 0;
        memory[ 6856] = 0;
        memory[ 6857] = 0;
        memory[ 6858] = 0;
        memory[ 6859] = 0;
        memory[ 6860] = 0;
        memory[ 6861] = 0;
        memory[ 6862] = 0;
        memory[ 6863] = 0;
        memory[ 6864] = 0;
        memory[ 6865] = 0;
        memory[ 6866] = 0;
        memory[ 6867] = 0;
        memory[ 6868] = 0;
        memory[ 6869] = 0;
        memory[ 6870] = 0;
        memory[ 6871] = 0;
        memory[ 6872] = 0;
        memory[ 6873] = 0;
        memory[ 6874] = 0;
        memory[ 6875] = 0;
        memory[ 6876] = 0;
        memory[ 6877] = 1;
        memory[ 6878] = 0;
        memory[ 6879] = 1;
        memory[ 6880] = 0;
        memory[ 6881] = 0;
        memory[ 6882] = 0;
        memory[ 6883] = 0;
        memory[ 6884] = 1;
        memory[ 6885] = 1;
        memory[ 6886] = 1;
        memory[ 6887] = 0;
        memory[ 6888] = 1;
        memory[ 6889] = 0;
        memory[ 6890] = 0;
        memory[ 6891] = 0;
        memory[ 6892] = 0;
        memory[ 6893] = 0;
        memory[ 6894] = 0;
        memory[ 6895] = 0;
        memory[ 6896] = 0;
        memory[ 6897] = 0;
        memory[ 6898] = 0;
        memory[ 6899] = 0;
        memory[ 6900] = 1;
        memory[ 6901] = 0;
        memory[ 6902] = 0;
        memory[ 6903] = 1;
        memory[ 6904] = 0;
        memory[ 6905] = 0;
        memory[ 6906] = 0;
        memory[ 6907] = 0;
        memory[ 6908] = 0;
        memory[ 6909] = 0;
        memory[ 6910] = 0;
        memory[ 6911] = 0;
        memory[ 6912] = 0;
        memory[ 6913] = 0;
        memory[ 6914] = 0;
        memory[ 6915] = 0;
        memory[ 6916] = 0;
        memory[ 6917] = 0;
        memory[ 6918] = 0;
        memory[ 6919] = 0;
        memory[ 6920] = 0;
        memory[ 6921] = 0;
        memory[ 6922] = 0;
        memory[ 6923] = 0;
        memory[ 6924] = 0;
        memory[ 6925] = 0;
        memory[ 6926] = 0;
        memory[ 6927] = 0;
        memory[ 6928] = 0;
        memory[ 6929] = 0;
        memory[ 6930] = 0;
        memory[ 6931] = 0;
        memory[ 6932] = 0;
        memory[ 6933] = 0;
        memory[ 6934] = 1;
        memory[ 6935] = 0;
        memory[ 6936] = 0;
        memory[ 6937] = 0;
        memory[ 6938] = 0;
        memory[ 6939] = 0;
        memory[ 6940] = 0;
        memory[ 6941] = 0;
        memory[ 6942] = 0;
        memory[ 6943] = 0;
        memory[ 6944] = 0;
        memory[ 6945] = 0;
        memory[ 6946] = 0;
        memory[ 6947] = 0;
        memory[ 6948] = 0;
        memory[ 6949] = 0;
        memory[ 6950] = 0;
        memory[ 6951] = 0;
        memory[ 6952] = 0;
        memory[ 6953] = 0;
        memory[ 6954] = 0;
        memory[ 6955] = 0;
        memory[ 6956] = 0;
        memory[ 6957] = 0;
        memory[ 6958] = 0;
        memory[ 6959] = 0;
        memory[ 6960] = 0;
        memory[ 6961] = 0;
        memory[ 6962] = 0;
        memory[ 6963] = 0;
        memory[ 6964] = 0;
        memory[ 6965] = 0;
        memory[ 6966] = 0;
        memory[ 6967] = 0;
        memory[ 6968] = 0;
        memory[ 6969] = 1;
        memory[ 6970] = 1;
        memory[ 6971] = 0;
        memory[ 6972] = 0;
        memory[ 6973] = 0;
        memory[ 6974] = 1;
        memory[ 6975] = 0;
        memory[ 6976] = 0;
        memory[ 6977] = 0;
        memory[ 6978] = 0;
        memory[ 6979] = 1;
        memory[ 6980] = 0;
        memory[ 6981] = 0;
        memory[ 6982] = 0;
        memory[ 6983] = 0;
        memory[ 6984] = 0;
        memory[ 6985] = 1;
        memory[ 6986] = 1;
        memory[ 6987] = 0;
        memory[ 6988] = 0;
        memory[ 6989] = 0;
        memory[ 6990] = 0;
        memory[ 6991] = 0;
        memory[ 6992] = 0;
        memory[ 6993] = 0;
        memory[ 6994] = 0;
        memory[ 6995] = 0;
        memory[ 6996] = 0;
        memory[ 6997] = 0;
        memory[ 6998] = 0;
        memory[ 6999] = 0;
        memory[ 7000] = 0;
        memory[ 7001] = 0;
        memory[ 7002] = 0;
        memory[ 7003] = 0;
        memory[ 7004] = 0;
        memory[ 7005] = 0;
        memory[ 7006] = 0;
        memory[ 7007] = 0;
        memory[ 7008] = 0;
        memory[ 7009] = 0;
        memory[ 7010] = 0;
        memory[ 7011] = 0;
        memory[ 7012] = 0;
        memory[ 7013] = 0;
        memory[ 7014] = 0;
        memory[ 7015] = 0;
        memory[ 7016] = 0;
        memory[ 7017] = 0;
        memory[ 7018] = 0;
        memory[ 7019] = 0;
        memory[ 7020] = 0;
        memory[ 7021] = 0;
        memory[ 7022] = 0;
        memory[ 7023] = 1;
        memory[ 7024] = 0;
        memory[ 7025] = 0;
        memory[ 7026] = 0;
        memory[ 7027] = 0;
        memory[ 7028] = 0;
        memory[ 7029] = 0;
        memory[ 7030] = 0;
        memory[ 7031] = 0;
        memory[ 7032] = 0;
        memory[ 7033] = 0;
        memory[ 7034] = 0;
        memory[ 7035] = 0;
        memory[ 7036] = 0;
        memory[ 7037] = 0;
        memory[ 7038] = 1;
        memory[ 7039] = 1;
        memory[ 7040] = 1;
        memory[ 7041] = 0;
        memory[ 7042] = 0;
        memory[ 7043] = 0;
        memory[ 7044] = 0;
        memory[ 7045] = 0;
        memory[ 7046] = 0;
        memory[ 7047] = 0;
        memory[ 7048] = 0;
        memory[ 7049] = 0;
        memory[ 7050] = 0;
        memory[ 7051] = 0;
        memory[ 7052] = 0;
        memory[ 7053] = 0;
        memory[ 7054] = 0;
        memory[ 7055] = 1;
        memory[ 7056] = 1;
        memory[ 7057] = 1;
        memory[ 7058] = 0;
        memory[ 7059] = 0;
        memory[ 7060] = 0;
        memory[ 7061] = 0;
        memory[ 7062] = 0;
        memory[ 7063] = 0;
        memory[ 7064] = 0;
        memory[ 7065] = 0;
        memory[ 7066] = 0;
        memory[ 7067] = 0;
        memory[ 7068] = 0;
        memory[ 7069] = 0;
        memory[ 7070] = 0;
        memory[ 7071] = 0;
        memory[ 7072] = 0;
        memory[ 7073] = 0;
        memory[ 7074] = 0;
        memory[ 7075] = 0;
        memory[ 7076] = 0;
        memory[ 7077] = 0;
        memory[ 7078] = 0;
        memory[ 7079] = 0;
        memory[ 7080] = 0;
        memory[ 7081] = 0;
        memory[ 7082] = 0;
        memory[ 7083] = 0;
        memory[ 7084] = 1;
        memory[ 7085] = 0;
        memory[ 7086] = 0;
        memory[ 7087] = 0;
        memory[ 7088] = 0;
        memory[ 7089] = 0;
        memory[ 7090] = 0;
        memory[ 7091] = 0;
        memory[ 7092] = 0;
        memory[ 7093] = 0;
        memory[ 7094] = 0;
        memory[ 7095] = 0;
        memory[ 7096] = 0;
        memory[ 7097] = 0;
        memory[ 7098] = 0;
        memory[ 7099] = 0;
        memory[ 7100] = 0;
        memory[ 7101] = 0;
        memory[ 7102] = 0;
        memory[ 7103] = 0;
        memory[ 7104] = 0;
        memory[ 7105] = 0;
        memory[ 7106] = 0;
        memory[ 7107] = 0;
        memory[ 7108] = 0;
        memory[ 7109] = 0;
        memory[ 7110] = 0;
        memory[ 7111] = 0;
        memory[ 7112] = 0;
        memory[ 7113] = 0;
        memory[ 7114] = 0;
        memory[ 7115] = 0;
        memory[ 7116] = 1;
        memory[ 7117] = 0;
        memory[ 7118] = 0;
        memory[ 7119] = 0;
        memory[ 7120] = 1;
        memory[ 7121] = 1;
        memory[ 7122] = 0;
        memory[ 7123] = 0;
        memory[ 7124] = 0;
        memory[ 7125] = 0;
        memory[ 7126] = 0;
        memory[ 7127] = 0;
        memory[ 7128] = 0;
        memory[ 7129] = 0;
        memory[ 7130] = 0;
        memory[ 7131] = 0;
        memory[ 7132] = 0;
        memory[ 7133] = 0;
        memory[ 7134] = 0;
        memory[ 7135] = 0;
        memory[ 7136] = 0;
        memory[ 7137] = 0;
        memory[ 7138] = 0;
        memory[ 7139] = 0;
        memory[ 7140] = 0;
        memory[ 7141] = 1;
        memory[ 7142] = 0;
        memory[ 7143] = 0;
        memory[ 7144] = 0;
        memory[ 7145] = 0;
        memory[ 7146] = 0;
        memory[ 7147] = 0;
        memory[ 7148] = 0;
        memory[ 7149] = 0;
        memory[ 7150] = 0;
        memory[ 7151] = 0;
        memory[ 7152] = 0;
        memory[ 7153] = 0;
        memory[ 7154] = 1;
        memory[ 7155] = 1;
        memory[ 7156] = 0;
        memory[ 7157] = 0;
        memory[ 7158] = 0;
        memory[ 7159] = 0;
        memory[ 7160] = 0;
        memory[ 7161] = 0;
        memory[ 7162] = 0;
        memory[ 7163] = 0;
        memory[ 7164] = 0;
        memory[ 7165] = 0;
        memory[ 7166] = 0;
        memory[ 7167] = 0;
        memory[ 7168] = 0;
        memory[ 7169] = 0;
        memory[ 7170] = 0;
        memory[ 7171] = 0;
        memory[ 7172] = 0;
        memory[ 7173] = 0;
        memory[ 7174] = 0;
        memory[ 7175] = 0;
        memory[ 7176] = 0;
        memory[ 7177] = 0;
        memory[ 7178] = 0;
        memory[ 7179] = 0;
        memory[ 7180] = 0;
        memory[ 7181] = 0;
        memory[ 7182] = 0;
        memory[ 7183] = 0;
        memory[ 7184] = 0;
        memory[ 7185] = 0;
        memory[ 7186] = 1;
        memory[ 7187] = 0;
        memory[ 7188] = 0;
        memory[ 7189] = 0;
        memory[ 7190] = 0;
        memory[ 7191] = 0;
        memory[ 7192] = 1;
        memory[ 7193] = 0;
        memory[ 7194] = 0;
        memory[ 7195] = 0;
        memory[ 7196] = 0;
        memory[ 7197] = 0;
        memory[ 7198] = 1;
        memory[ 7199] = 1;
        memory[ 7200] = 0;
        memory[ 7201] = 0;
        memory[ 7202] = 0;
        memory[ 7203] = 1;
        memory[ 7204] = 1;
        memory[ 7205] = 0;
        memory[ 7206] = 1;
        memory[ 7207] = 1;
        memory[ 7208] = 0;
        memory[ 7209] = 0;
        memory[ 7210] = 0;
        memory[ 7211] = 1;
        memory[ 7212] = 0;
        memory[ 7213] = 0;
        memory[ 7214] = 0;
        memory[ 7215] = 0;
        memory[ 7216] = 0;
        memory[ 7217] = 0;
        memory[ 7218] = 0;
        memory[ 7219] = 0;
        memory[ 7220] = 0;
        memory[ 7221] = 0;
        memory[ 7222] = 0;
        memory[ 7223] = 0;
        memory[ 7224] = 0;
        memory[ 7225] = 0;
        memory[ 7226] = 0;
        memory[ 7227] = 1;
        memory[ 7228] = 0;
        memory[ 7229] = 0;
        memory[ 7230] = 0;
        memory[ 7231] = 0;
        memory[ 7232] = 0;
        memory[ 7233] = 1;
        memory[ 7234] = 0;
        memory[ 7235] = 0;
        memory[ 7236] = 0;
        memory[ 7237] = 0;
        memory[ 7238] = 0;
        memory[ 7239] = 0;
        memory[ 7240] = 0;
        memory[ 7241] = 0;
        memory[ 7242] = 0;
        memory[ 7243] = 1;
        memory[ 7244] = 1;
        memory[ 7245] = 0;
        memory[ 7246] = 0;
        memory[ 7247] = 0;
        memory[ 7248] = 0;
        memory[ 7249] = 0;
        memory[ 7250] = 0;
        memory[ 7251] = 0;
        memory[ 7252] = 0;
        memory[ 7253] = 0;
        memory[ 7254] = 0;
        memory[ 7255] = 1;
        memory[ 7256] = 1;
        memory[ 7257] = 1;
        memory[ 7258] = 0;
        memory[ 7259] = 0;
        memory[ 7260] = 0;
        memory[ 7261] = 0;
        memory[ 7262] = 0;
        memory[ 7263] = 0;
        memory[ 7264] = 0;
        memory[ 7265] = 0;
        memory[ 7266] = 0;
        memory[ 7267] = 0;
        memory[ 7268] = 0;
        memory[ 7269] = 0;
        memory[ 7270] = 0;
        memory[ 7271] = 0;
        memory[ 7272] = 0;
        memory[ 7273] = 0;
        memory[ 7274] = 0;
        memory[ 7275] = 0;
        memory[ 7276] = 0;
        memory[ 7277] = 0;
        memory[ 7278] = 0;
        memory[ 7279] = 1;
        memory[ 7280] = 0;
        memory[ 7281] = 0;
        memory[ 7282] = 0;
        memory[ 7283] = 0;
        memory[ 7284] = 1;
        memory[ 7285] = 1;
        memory[ 7286] = 0;
        memory[ 7287] = 0;
        memory[ 7288] = 0;
        memory[ 7289] = 0;
        memory[ 7290] = 0;
        memory[ 7291] = 1;
        memory[ 7292] = 0;
        memory[ 7293] = 0;
        memory[ 7294] = 0;
        memory[ 7295] = 0;
        memory[ 7296] = 0;
        memory[ 7297] = 0;
        memory[ 7298] = 0;
        memory[ 7299] = 0;
        memory[ 7300] = 0;
        memory[ 7301] = 0;
        memory[ 7302] = 0;
        memory[ 7303] = 0;
        memory[ 7304] = 0;
        memory[ 7305] = 1;
        memory[ 7306] = 0;
        memory[ 7307] = 0;
        memory[ 7308] = 0;
        memory[ 7309] = 0;
        memory[ 7310] = 0;
        memory[ 7311] = 0;
        memory[ 7312] = 0;
        memory[ 7313] = 1;
        memory[ 7314] = 0;
        memory[ 7315] = 0;
        memory[ 7316] = 0;
        memory[ 7317] = 0;
        memory[ 7318] = 0;
        memory[ 7319] = 0;
        memory[ 7320] = 0;
        memory[ 7321] = 0;
        memory[ 7322] = 0;
        memory[ 7323] = 0;
        memory[ 7324] = 0;
        memory[ 7325] = 0;
        memory[ 7326] = 0;
        memory[ 7327] = 0;
        memory[ 7328] = 0;
        memory[ 7329] = 0;
        memory[ 7330] = 0;
        memory[ 7331] = 0;
        memory[ 7332] = 0;
        memory[ 7333] = 0;
        memory[ 7334] = 0;
        memory[ 7335] = 0;
        memory[ 7336] = 0;
        memory[ 7337] = 0;
        memory[ 7338] = 1;
        memory[ 7339] = 0;
        memory[ 7340] = 0;
        memory[ 7341] = 0;
        memory[ 7342] = 0;
        memory[ 7343] = 0;
        memory[ 7344] = 0;
        memory[ 7345] = 0;
        memory[ 7346] = 0;
        memory[ 7347] = 0;
        memory[ 7348] = 0;
        memory[ 7349] = 0;
        memory[ 7350] = 0;
        memory[ 7351] = 0;
        memory[ 7352] = 0;
        memory[ 7353] = 0;
        memory[ 7354] = 0;
        memory[ 7355] = 0;
        memory[ 7356] = 0;
        memory[ 7357] = 0;
        memory[ 7358] = 0;
        memory[ 7359] = 0;
        memory[ 7360] = 0;
        memory[ 7361] = 0;
        memory[ 7362] = 0;
        memory[ 7363] = 0;
        memory[ 7364] = 0;
        memory[ 7365] = 0;
        memory[ 7366] = 0;
        memory[ 7367] = 0;
        memory[ 7368] = 0;
        memory[ 7369] = 1;
        memory[ 7370] = 1;
        memory[ 7371] = 0;
        memory[ 7372] = 0;
        memory[ 7373] = 0;
        memory[ 7374] = 0;
        memory[ 7375] = 0;
        memory[ 7376] = 1;
        memory[ 7377] = 1;
        memory[ 7378] = 0;
        memory[ 7379] = 0;
        memory[ 7380] = 0;
        memory[ 7381] = 0;
        memory[ 7382] = 0;
        memory[ 7383] = 0;
        memory[ 7384] = 0;
        memory[ 7385] = 0;
        memory[ 7386] = 0;
        memory[ 7387] = 0;
        memory[ 7388] = 0;
        memory[ 7389] = 0;
        memory[ 7390] = 0;
        memory[ 7391] = 0;
        memory[ 7392] = 0;
        memory[ 7393] = 0;
        memory[ 7394] = 0;
        memory[ 7395] = 0;
        memory[ 7396] = 0;
        memory[ 7397] = 0;
        memory[ 7398] = 0;
        memory[ 7399] = 0;
        memory[ 7400] = 1;
        memory[ 7401] = 0;
        memory[ 7402] = 0;
        memory[ 7403] = 0;
        memory[ 7404] = 0;
        memory[ 7405] = 1;
        memory[ 7406] = 0;
        memory[ 7407] = 0;
        memory[ 7408] = 1;
        memory[ 7409] = 0;
        memory[ 7410] = 0;
        memory[ 7411] = 0;
        memory[ 7412] = 0;
        memory[ 7413] = 0;
        memory[ 7414] = 0;
        memory[ 7415] = 0;
        memory[ 7416] = 0;
        memory[ 7417] = 0;
        memory[ 7418] = 0;
        memory[ 7419] = 1;
        memory[ 7420] = 0;
        memory[ 7421] = 0;
        memory[ 7422] = 1;
        memory[ 7423] = 0;
        memory[ 7424] = 0;
        memory[ 7425] = 0;
        memory[ 7426] = 0;
        memory[ 7427] = 0;
        memory[ 7428] = 0;
        memory[ 7429] = 0;
        memory[ 7430] = 0;
        memory[ 7431] = 1;
        memory[ 7432] = 0;
        memory[ 7433] = 0;
        memory[ 7434] = 0;
        memory[ 7435] = 0;
        memory[ 7436] = 0;
        memory[ 7437] = 0;
        memory[ 7438] = 0;
        memory[ 7439] = 0;
        memory[ 7440] = 0;
        memory[ 7441] = 0;
        memory[ 7442] = 0;
        memory[ 7443] = 0;
        memory[ 7444] = 0;
        memory[ 7445] = 0;
        memory[ 7446] = 0;
        memory[ 7447] = 0;
        memory[ 7448] = 0;
        memory[ 7449] = 0;
        memory[ 7450] = 0;
        memory[ 7451] = 0;
        memory[ 7452] = 0;
        memory[ 7453] = 0;
        memory[ 7454] = 0;
        memory[ 7455] = 0;
        memory[ 7456] = 0;
        memory[ 7457] = 0;
        memory[ 7458] = 0;
        memory[ 7459] = 0;
        memory[ 7460] = 0;
        memory[ 7461] = 0;
        memory[ 7462] = 0;
        memory[ 7463] = 0;
        memory[ 7464] = 0;
        memory[ 7465] = 0;
        memory[ 7466] = 0;
        memory[ 7467] = 0;
        memory[ 7468] = 0;
        memory[ 7469] = 1;
        memory[ 7470] = 0;
        memory[ 7471] = 0;
        memory[ 7472] = 0;
        memory[ 7473] = 0;
        memory[ 7474] = 0;
        memory[ 7475] = 0;
        memory[ 7476] = 0;
        memory[ 7477] = 0;
        memory[ 7478] = 0;
        memory[ 7479] = 0;
        memory[ 7480] = 0;
        memory[ 7481] = 0;
        memory[ 7482] = 0;
        memory[ 7483] = 0;
        memory[ 7484] = 0;
        memory[ 7485] = 0;
        memory[ 7486] = 1;
        memory[ 7487] = 0;
        memory[ 7488] = 0;
        memory[ 7489] = 0;
        memory[ 7490] = 0;
        memory[ 7491] = 0;
        memory[ 7492] = 0;
        memory[ 7493] = 0;
        memory[ 7494] = 0;
        memory[ 7495] = 0;
        memory[ 7496] = 0;
        memory[ 7497] = 0;
        memory[ 7498] = 0;
        memory[ 7499] = 0;
        memory[ 7500] = 0;
        memory[ 7501] = 0;
        memory[ 7502] = 0;
        memory[ 7503] = 0;
        memory[ 7504] = 0;
        memory[ 7505] = 0;
        memory[ 7506] = 0;
        memory[ 7507] = 0;
        memory[ 7508] = 0;
        memory[ 7509] = 0;
        memory[ 7510] = 0;
        memory[ 7511] = 0;
        memory[ 7512] = 0;
        memory[ 7513] = 1;
        memory[ 7514] = 1;
        memory[ 7515] = 1;
        memory[ 7516] = 0;
        memory[ 7517] = 1;
        memory[ 7518] = 1;
        memory[ 7519] = 1;
        memory[ 7520] = 0;
        memory[ 7521] = 0;
        memory[ 7522] = 0;
        memory[ 7523] = 0;
        memory[ 7524] = 0;
        memory[ 7525] = 0;
        memory[ 7526] = 0;
        memory[ 7527] = 0;
        memory[ 7528] = 1;
        memory[ 7529] = 0;
        memory[ 7530] = 0;
        memory[ 7531] = 0;
        memory[ 7532] = 0;
        memory[ 7533] = 0;
        memory[ 7534] = 0;
        memory[ 7535] = 1;
        memory[ 7536] = 0;
        memory[ 7537] = 0;
        memory[ 7538] = 0;
        memory[ 7539] = 0;
        memory[ 7540] = 0;
        memory[ 7541] = 0;
        memory[ 7542] = 0;
        memory[ 7543] = 0;
        memory[ 7544] = 0;
        memory[ 7545] = 0;
        memory[ 7546] = 0;
        memory[ 7547] = 0;
        memory[ 7548] = 0;
        memory[ 7549] = 0;
        memory[ 7550] = 0;
        memory[ 7551] = 0;
        memory[ 7552] = 0;
        memory[ 7553] = 0;
        memory[ 7554] = 0;
        memory[ 7555] = 0;
        memory[ 7556] = 0;
        memory[ 7557] = 0;
        memory[ 7558] = 0;
        memory[ 7559] = 0;
        memory[ 7560] = 0;
        memory[ 7561] = 0;
        memory[ 7562] = 0;
        memory[ 7563] = 0;
        memory[ 7564] = 0;
        memory[ 7565] = 0;
        memory[ 7566] = 0;
        memory[ 7567] = 0;
        memory[ 7568] = 0;
        memory[ 7569] = 0;
        memory[ 7570] = 0;
        memory[ 7571] = 0;
        memory[ 7572] = 0;
        memory[ 7573] = 0;
        memory[ 7574] = 0;
        memory[ 7575] = 1;
        memory[ 7576] = 1;
        memory[ 7577] = 0;
        memory[ 7578] = 0;
        memory[ 7579] = 0;
        memory[ 7580] = 1;
        memory[ 7581] = 1;
        memory[ 7582] = 0;
        memory[ 7583] = 0;
        memory[ 7584] = 0;
        memory[ 7585] = 0;
        memory[ 7586] = 0;
        memory[ 7587] = 0;
        memory[ 7588] = 0;
        memory[ 7589] = 0;
        memory[ 7590] = 1;
        memory[ 7591] = 0;
        memory[ 7592] = 0;
        memory[ 7593] = 0;
        memory[ 7594] = 0;
        memory[ 7595] = 0;
        memory[ 7596] = 0;
        memory[ 7597] = 0;
        memory[ 7598] = 0;
        memory[ 7599] = 0;
        memory[ 7600] = 0;
        memory[ 7601] = 0;
        memory[ 7602] = 0;
        memory[ 7603] = 0;
        memory[ 7604] = 1;
        memory[ 7605] = 1;
        memory[ 7606] = 1;
        memory[ 7607] = 1;
        memory[ 7608] = 0;
        memory[ 7609] = 0;
        memory[ 7610] = 0;
        memory[ 7611] = 0;
        memory[ 7612] = 1;
        memory[ 7613] = 0;
        memory[ 7614] = 0;
        memory[ 7615] = 0;
        memory[ 7616] = 0;
        memory[ 7617] = 0;
        memory[ 7618] = 0;
        memory[ 7619] = 0;
        memory[ 7620] = 0;
        memory[ 7621] = 0;
        memory[ 7622] = 0;
        memory[ 7623] = 0;
        memory[ 7624] = 0;
        memory[ 7625] = 0;
        memory[ 7626] = 0;
        memory[ 7627] = 0;
        memory[ 7628] = 0;
        memory[ 7629] = 0;
        memory[ 7630] = 0;
        memory[ 7631] = 0;
        memory[ 7632] = 0;
        memory[ 7633] = 0;
        memory[ 7634] = 0;
        memory[ 7635] = 0;
        memory[ 7636] = 1;
        memory[ 7637] = 0;
        memory[ 7638] = 1;
        memory[ 7639] = 0;
        memory[ 7640] = 0;
        memory[ 7641] = 0;
        memory[ 7642] = 0;
        memory[ 7643] = 0;
        memory[ 7644] = 0;
        memory[ 7645] = 0;
        memory[ 7646] = 0;
        memory[ 7647] = 0;
        memory[ 7648] = 1;
        memory[ 7649] = 1;
        memory[ 7650] = 0;
        memory[ 7651] = 0;
        memory[ 7652] = 0;
        memory[ 7653] = 0;
        memory[ 7654] = 0;
        memory[ 7655] = 0;
        memory[ 7656] = 0;
        memory[ 7657] = 0;
        memory[ 7658] = 0;
        memory[ 7659] = 0;
        memory[ 7660] = 0;
        memory[ 7661] = 1;
        memory[ 7662] = 0;
        memory[ 7663] = 1;
        memory[ 7664] = 0;
        memory[ 7665] = 1;
        memory[ 7666] = 1;
        memory[ 7667] = 1;
        memory[ 7668] = 1;
        memory[ 7669] = 0;
        memory[ 7670] = 0;
        memory[ 7671] = 0;
        memory[ 7672] = 0;
        memory[ 7673] = 0;
        memory[ 7674] = 0;
        memory[ 7675] = 1;
        memory[ 7676] = 0;
        memory[ 7677] = 0;
        memory[ 7678] = 0;
        memory[ 7679] = 0;
        memory[ 7680] = 0;
        memory[ 7681] = 0;
        memory[ 7682] = 0;
        memory[ 7683] = 0;
        memory[ 7684] = 0;
        memory[ 7685] = 0;
        memory[ 7686] = 0;
        memory[ 7687] = 0;
        memory[ 7688] = 1;
        memory[ 7689] = 0;
        memory[ 7690] = 0;
        memory[ 7691] = 1;
        memory[ 7692] = 0;
        memory[ 7693] = 1;
        memory[ 7694] = 1;
        memory[ 7695] = 0;
        memory[ 7696] = 0;
        memory[ 7697] = 0;
        memory[ 7698] = 0;
        memory[ 7699] = 0;
        memory[ 7700] = 0;
        memory[ 7701] = 0;
        memory[ 7702] = 0;
        memory[ 7703] = 0;
        memory[ 7704] = 0;
        memory[ 7705] = 0;
        memory[ 7706] = 0;
        memory[ 7707] = 0;
        memory[ 7708] = 0;
        memory[ 7709] = 0;
        memory[ 7710] = 0;
        memory[ 7711] = 0;
        memory[ 7712] = 0;
        memory[ 7713] = 0;
        memory[ 7714] = 0;
        memory[ 7715] = 0;
        memory[ 7716] = 0;
        memory[ 7717] = 0;
        memory[ 7718] = 0;
        memory[ 7719] = 0;
        memory[ 7720] = 0;
        memory[ 7721] = 0;
        memory[ 7722] = 0;
        memory[ 7723] = 0;
        memory[ 7724] = 0;
        memory[ 7725] = 0;
        memory[ 7726] = 0;
        memory[ 7727] = 0;
        memory[ 7728] = 0;
        memory[ 7729] = 1;
        memory[ 7730] = 0;
        memory[ 7731] = 0;
        memory[ 7732] = 1;
        memory[ 7733] = 0;
        memory[ 7734] = 0;
        memory[ 7735] = 0;
        memory[ 7736] = 0;
        memory[ 7737] = 0;
        memory[ 7738] = 0;
        memory[ 7739] = 0;
        memory[ 7740] = 0;
        memory[ 7741] = 1;
        memory[ 7742] = 0;
        memory[ 7743] = 0;
        memory[ 7744] = 0;
        memory[ 7745] = 0;
        memory[ 7746] = 0;
        memory[ 7747] = 0;
        memory[ 7748] = 0;
        memory[ 7749] = 0;
        memory[ 7750] = 0;
        memory[ 7751] = 0;
        memory[ 7752] = 0;
        memory[ 7753] = 0;
        memory[ 7754] = 0;
        memory[ 7755] = 0;
        memory[ 7756] = 0;
        memory[ 7757] = 1;
        memory[ 7758] = 0;
        memory[ 7759] = 0;
        memory[ 7760] = 0;
        memory[ 7761] = 0;
        memory[ 7762] = 1;
        memory[ 7763] = 0;
        memory[ 7764] = 0;
        memory[ 7765] = 0;
        memory[ 7766] = 1;
        memory[ 7767] = 0;
        memory[ 7768] = 0;
        memory[ 7769] = 0;
        memory[ 7770] = 1;
        memory[ 7771] = 0;
        memory[ 7772] = 0;
        memory[ 7773] = 0;
        memory[ 7774] = 0;
        memory[ 7775] = 0;
        memory[ 7776] = 0;
        memory[ 7777] = 0;
        memory[ 7778] = 0;
        memory[ 7779] = 0;
        memory[ 7780] = 0;
        memory[ 7781] = 0;
        memory[ 7782] = 0;
        memory[ 7783] = 0;
        memory[ 7784] = 0;
        memory[ 7785] = 0;
        memory[ 7786] = 0;
        memory[ 7787] = 1;
        memory[ 7788] = 0;
        memory[ 7789] = 0;
        memory[ 7790] = 0;
        memory[ 7791] = 0;
        memory[ 7792] = 0;
        memory[ 7793] = 0;
        memory[ 7794] = 0;
        memory[ 7795] = 0;
        memory[ 7796] = 0;
        memory[ 7797] = 0;
        memory[ 7798] = 0;
        memory[ 7799] = 0;
        memory[ 7800] = 0;
        memory[ 7801] = 0;
        memory[ 7802] = 0;
        memory[ 7803] = 0;
        memory[ 7804] = 0;
        memory[ 7805] = 0;
        memory[ 7806] = 0;
        memory[ 7807] = 0;
        memory[ 7808] = 0;
        memory[ 7809] = 0;
        memory[ 7810] = 0;
        memory[ 7811] = 0;
        memory[ 7812] = 0;
        memory[ 7813] = 0;
        memory[ 7814] = 0;
        memory[ 7815] = 0;
        memory[ 7816] = 0;
        memory[ 7817] = 0;
        memory[ 7818] = 0;
        memory[ 7819] = 0;
        memory[ 7820] = 0;
        memory[ 7821] = 0;
        memory[ 7822] = 0;
        memory[ 7823] = 0;
        memory[ 7824] = 0;
        memory[ 7825] = 0;
        memory[ 7826] = 0;
        memory[ 7827] = 0;
        memory[ 7828] = 0;
        memory[ 7829] = 0;
        memory[ 7830] = 0;
        memory[ 7831] = 1;
        memory[ 7832] = 0;
        memory[ 7833] = 0;
        memory[ 7834] = 0;
        memory[ 7835] = 0;
        memory[ 7836] = 0;
        memory[ 7837] = 0;
        memory[ 7838] = 0;
        memory[ 7839] = 0;
        memory[ 7840] = 0;
        memory[ 7841] = 0;
        memory[ 7842] = 0;
        memory[ 7843] = 0;
        memory[ 7844] = 0;
        memory[ 7845] = 0;
        memory[ 7846] = 0;
        memory[ 7847] = 0;
        memory[ 7848] = 0;
        memory[ 7849] = 0;
        memory[ 7850] = 0;
        memory[ 7851] = 0;
        memory[ 7852] = 0;
        memory[ 7853] = 1;
        memory[ 7854] = 1;
        memory[ 7855] = 0;
        memory[ 7856] = 0;
        memory[ 7857] = 0;
        memory[ 7858] = 0;
        memory[ 7859] = 0;
        memory[ 7860] = 1;
        memory[ 7861] = 0;
        memory[ 7862] = 0;
        memory[ 7863] = 0;
        memory[ 7864] = 0;
        memory[ 7865] = 0;
        memory[ 7866] = 0;
        memory[ 7867] = 0;
        memory[ 7868] = 1;
        memory[ 7869] = 0;
        memory[ 7870] = 0;
        memory[ 7871] = 0;
        memory[ 7872] = 0;
        memory[ 7873] = 0;
        memory[ 7874] = 0;
        memory[ 7875] = 0;
        memory[ 7876] = 0;
        memory[ 7877] = 0;
        memory[ 7878] = 0;
        memory[ 7879] = 0;
        memory[ 7880] = 0;
        memory[ 7881] = 0;
        memory[ 7882] = 0;
        memory[ 7883] = 0;
        memory[ 7884] = 0;
        memory[ 7885] = 0;
        memory[ 7886] = 0;
        memory[ 7887] = 0;
        memory[ 7888] = 0;
        memory[ 7889] = 0;
        memory[ 7890] = 0;
        memory[ 7891] = 0;
        memory[ 7892] = 0;
        memory[ 7893] = 0;
        memory[ 7894] = 0;
        memory[ 7895] = 0;
        memory[ 7896] = 0;
        memory[ 7897] = 0;
        memory[ 7898] = 0;
        memory[ 7899] = 0;
        memory[ 7900] = 0;
        memory[ 7901] = 0;
        memory[ 7902] = 0;
        memory[ 7903] = 0;
        memory[ 7904] = 0;
        memory[ 7905] = 0;
        memory[ 7906] = 0;
        memory[ 7907] = 0;
        memory[ 7908] = 0;
        memory[ 7909] = 0;
        memory[ 7910] = 0;
        memory[ 7911] = 0;
        memory[ 7912] = 0;
        memory[ 7913] = 0;
        memory[ 7914] = 0;
        memory[ 7915] = 0;
        memory[ 7916] = 0;
        memory[ 7917] = 1;
        memory[ 7918] = 0;
        memory[ 7919] = 0;
        memory[ 7920] = 0;
        memory[ 7921] = 1;
        memory[ 7922] = 0;
        memory[ 7923] = 0;
        memory[ 7924] = 0;
        memory[ 7925] = 0;
        memory[ 7926] = 0;
        memory[ 7927] = 0;
        memory[ 7928] = 0;
        memory[ 7929] = 0;
        memory[ 7930] = 0;
        memory[ 7931] = 0;
        memory[ 7932] = 0;
        memory[ 7933] = 0;
        memory[ 7934] = 0;
        memory[ 7935] = 0;
        memory[ 7936] = 0;
        memory[ 7937] = 0;
        memory[ 7938] = 0;
        memory[ 7939] = 0;
        memory[ 7940] = 0;
        memory[ 7941] = 0;
        memory[ 7942] = 0;
        memory[ 7943] = 0;
        memory[ 7944] = 0;
        memory[ 7945] = 0;
        memory[ 7946] = 0;
        memory[ 7947] = 0;
        memory[ 7948] = 0;
        memory[ 7949] = 1;
        memory[ 7950] = 1;
        memory[ 7951] = 0;
        memory[ 7952] = 0;
        memory[ 7953] = 0;
        memory[ 7954] = 0;
        memory[ 7955] = 0;
        memory[ 7956] = 0;
        memory[ 7957] = 1;
        memory[ 7958] = 1;
        memory[ 7959] = 0;
        memory[ 7960] = 0;
        memory[ 7961] = 0;
        memory[ 7962] = 0;
        memory[ 7963] = 0;
        memory[ 7964] = 0;
        memory[ 7965] = 0;
        memory[ 7966] = 0;
        memory[ 7967] = 0;
        memory[ 7968] = 0;
        memory[ 7969] = 0;
        memory[ 7970] = 0;
        memory[ 7971] = 0;
        memory[ 7972] = 0;
        memory[ 7973] = 0;
        memory[ 7974] = 0;
        memory[ 7975] = 0;
        memory[ 7976] = 0;
        memory[ 7977] = 0;
        memory[ 7978] = 1;
        memory[ 7979] = 1;
        memory[ 7980] = 0;
        memory[ 7981] = 0;
        memory[ 7982] = 0;
        memory[ 7983] = 0;
        memory[ 7984] = 0;
        memory[ 7985] = 0;
        memory[ 7986] = 1;
        memory[ 7987] = 1;
        memory[ 7988] = 1;
        memory[ 7989] = 0;
        memory[ 7990] = 0;
        memory[ 7991] = 1;
        memory[ 7992] = 0;
        memory[ 7993] = 0;
        memory[ 7994] = 0;
        memory[ 7995] = 0;
        memory[ 7996] = 0;
        memory[ 7997] = 0;
        memory[ 7998] = 0;
        memory[ 7999] = 0;
        memory[ 8000] = 0;
        memory[ 8001] = 0;
        memory[ 8002] = 0;
        memory[ 8003] = 0;
        memory[ 8004] = 1;
        memory[ 8005] = 0;
        memory[ 8006] = 0;
        memory[ 8007] = 0;
        memory[ 8008] = 0;
        memory[ 8009] = 1;
        memory[ 8010] = 1;
        memory[ 8011] = 0;
        memory[ 8012] = 0;
        memory[ 8013] = 0;
        memory[ 8014] = 0;
        memory[ 8015] = 0;
        memory[ 8016] = 0;
        memory[ 8017] = 0;
        memory[ 8018] = 0;
        memory[ 8019] = 0;
        memory[ 8020] = 0;
        memory[ 8021] = 0;
        memory[ 8022] = 0;
        memory[ 8023] = 0;
        memory[ 8024] = 0;
        memory[ 8025] = 0;
        memory[ 8026] = 0;
        memory[ 8027] = 0;
        memory[ 8028] = 0;
        memory[ 8029] = 0;
        memory[ 8030] = 0;
        memory[ 8031] = 0;
        memory[ 8032] = 0;
        memory[ 8033] = 0;
        memory[ 8034] = 0;
        memory[ 8035] = 0;
        memory[ 8036] = 0;
        memory[ 8037] = 1;
        memory[ 8038] = 0;
        memory[ 8039] = 1;
        memory[ 8040] = 1;
        memory[ 8041] = 1;
        memory[ 8042] = 0;
        memory[ 8043] = 0;
        memory[ 8044] = 0;
        memory[ 8045] = 0;
        memory[ 8046] = 0;
        memory[ 8047] = 0;
        memory[ 8048] = 0;
        memory[ 8049] = 0;
        memory[ 8050] = 0;
        memory[ 8051] = 0;
        memory[ 8052] = 0;
        memory[ 8053] = 0;
        memory[ 8054] = 0;
        memory[ 8055] = 0;
        memory[ 8056] = 0;
        memory[ 8057] = 0;
        memory[ 8058] = 0;
        memory[ 8059] = 1;
        memory[ 8060] = 1;
        memory[ 8061] = 0;
        memory[ 8062] = 0;
        memory[ 8063] = 0;
        memory[ 8064] = 0;
        memory[ 8065] = 0;
        memory[ 8066] = 0;
        memory[ 8067] = 0;
        memory[ 8068] = 0;
        memory[ 8069] = 0;
        memory[ 8070] = 0;
        memory[ 8071] = 0;
        memory[ 8072] = 0;
        memory[ 8073] = 0;
        memory[ 8074] = 0;
        memory[ 8075] = 0;
        memory[ 8076] = 0;
        memory[ 8077] = 0;
        memory[ 8078] = 0;
        memory[ 8079] = 0;
        memory[ 8080] = 0;
        memory[ 8081] = 1;
        memory[ 8082] = 0;
        memory[ 8083] = 0;
        memory[ 8084] = 0;
        memory[ 8085] = 0;
        memory[ 8086] = 0;
        memory[ 8087] = 1;
        memory[ 8088] = 0;
        memory[ 8089] = 0;
        memory[ 8090] = 0;
        memory[ 8091] = 0;
        memory[ 8092] = 0;
        memory[ 8093] = 0;
        memory[ 8094] = 0;
        memory[ 8095] = 0;
        memory[ 8096] = 0;
        memory[ 8097] = 0;
        memory[ 8098] = 0;
        memory[ 8099] = 0;
        memory[ 8100] = 0;
        memory[ 8101] = 1;
        memory[ 8102] = 0;
        memory[ 8103] = 0;
        memory[ 8104] = 0;
        memory[ 8105] = 0;
        memory[ 8106] = 0;
        memory[ 8107] = 0;
        memory[ 8108] = 0;
        memory[ 8109] = 0;
        memory[ 8110] = 1;
        memory[ 8111] = 1;
        memory[ 8112] = 0;
        memory[ 8113] = 0;
        memory[ 8114] = 0;
        memory[ 8115] = 1;
        memory[ 8116] = 1;
        memory[ 8117] = 0;
        memory[ 8118] = 0;
        memory[ 8119] = 1;
        memory[ 8120] = 0;
        memory[ 8121] = 0;
        memory[ 8122] = 0;
        memory[ 8123] = 0;
        memory[ 8124] = 0;
        memory[ 8125] = 0;
        memory[ 8126] = 0;
        memory[ 8127] = 0;
        memory[ 8128] = 0;
        memory[ 8129] = 0;
        memory[ 8130] = 0;
        memory[ 8131] = 0;
        memory[ 8132] = 0;
        memory[ 8133] = 0;
        memory[ 8134] = 0;
        memory[ 8135] = 0;
        memory[ 8136] = 0;
        memory[ 8137] = 0;
        memory[ 8138] = 1;
        memory[ 8139] = 0;
        memory[ 8140] = 0;
        memory[ 8141] = 0;
        memory[ 8142] = 0;
        memory[ 8143] = 0;
        memory[ 8144] = 0;
        memory[ 8145] = 0;
        memory[ 8146] = 0;
        memory[ 8147] = 0;
        memory[ 8148] = 0;
        memory[ 8149] = 0;
        memory[ 8150] = 0;
        memory[ 8151] = 0;
        memory[ 8152] = 0;
        memory[ 8153] = 0;
        memory[ 8154] = 1;
        memory[ 8155] = 0;
        memory[ 8156] = 0;
        memory[ 8157] = 0;
        memory[ 8158] = 1;
        memory[ 8159] = 1;
        memory[ 8160] = 1;
        memory[ 8161] = 0;
        memory[ 8162] = 0;
        memory[ 8163] = 0;
        memory[ 8164] = 0;
        memory[ 8165] = 0;
        memory[ 8166] = 0;
        memory[ 8167] = 0;
        memory[ 8168] = 0;
        memory[ 8169] = 0;
        memory[ 8170] = 0;
        memory[ 8171] = 0;
        memory[ 8172] = 0;
        memory[ 8173] = 0;
        memory[ 8174] = 0;
        memory[ 8175] = 0;
        memory[ 8176] = 0;
        memory[ 8177] = 0;
        memory[ 8178] = 0;
        memory[ 8179] = 0;
        memory[ 8180] = 0;
        memory[ 8181] = 0;
        memory[ 8182] = 0;
        memory[ 8183] = 0;
        memory[ 8184] = 0;
        memory[ 8185] = 0;
        memory[ 8186] = 0;
        memory[ 8187] = 0;
        memory[ 8188] = 1;
        memory[ 8189] = 0;
        memory[ 8190] = 0;
        memory[ 8191] = 0;
        memory[ 8192] = 0;
        memory[ 8193] = 0;
        memory[ 8194] = 0;
        memory[ 8195] = 0;
        memory[ 8196] = 1;
        memory[ 8197] = 0;
        memory[ 8198] = 1;
        memory[ 8199] = 0;
        memory[ 8200] = 0;
        memory[ 8201] = 0;
        memory[ 8202] = 0;
        memory[ 8203] = 0;
        memory[ 8204] = 0;
        memory[ 8205] = 0;
        memory[ 8206] = 0;
        memory[ 8207] = 0;
        memory[ 8208] = 0;
        memory[ 8209] = 1;
        memory[ 8210] = 0;
        memory[ 8211] = 0;
        memory[ 8212] = 0;
        memory[ 8213] = 0;
        memory[ 8214] = 0;
        memory[ 8215] = 0;
        memory[ 8216] = 0;
        memory[ 8217] = 1;
        memory[ 8218] = 1;
        memory[ 8219] = 0;
        memory[ 8220] = 1;
        memory[ 8221] = 0;
        memory[ 8222] = 0;
        memory[ 8223] = 0;
        memory[ 8224] = 0;
        memory[ 8225] = 0;
        memory[ 8226] = 0;
        memory[ 8227] = 0;
        memory[ 8228] = 0;
        memory[ 8229] = 0;
        memory[ 8230] = 0;
        memory[ 8231] = 0;
        memory[ 8232] = 0;
        memory[ 8233] = 0;
        memory[ 8234] = 0;
        memory[ 8235] = 0;
        memory[ 8236] = 0;
        memory[ 8237] = 0;
        memory[ 8238] = 1;
        memory[ 8239] = 0;
        memory[ 8240] = 0;
        memory[ 8241] = 0;
        memory[ 8242] = 0;
        memory[ 8243] = 0;
        memory[ 8244] = 0;
        memory[ 8245] = 0;
        memory[ 8246] = 0;
        memory[ 8247] = 0;
        memory[ 8248] = 0;
        memory[ 8249] = 0;
        memory[ 8250] = 0;
        memory[ 8251] = 0;
        memory[ 8252] = 0;
        memory[ 8253] = 0;
        memory[ 8254] = 0;
        memory[ 8255] = 0;
        memory[ 8256] = 0;
        memory[ 8257] = 0;
        memory[ 8258] = 0;
        memory[ 8259] = 0;
        memory[ 8260] = 0;
        memory[ 8261] = 0;
        memory[ 8262] = 0;
        memory[ 8263] = 0;
        memory[ 8264] = 0;
        memory[ 8265] = 0;
        memory[ 8266] = 0;
        memory[ 8267] = 0;
        memory[ 8268] = 0;
        memory[ 8269] = 0;
        memory[ 8270] = 0;
        memory[ 8271] = 0;
        memory[ 8272] = 0;
        memory[ 8273] = 0;
        memory[ 8274] = 0;
        memory[ 8275] = 0;
        memory[ 8276] = 0;
        memory[ 8277] = 0;
        memory[ 8278] = 0;
        memory[ 8279] = 0;
        memory[ 8280] = 0;
        memory[ 8281] = 0;
        memory[ 8282] = 0;
        memory[ 8283] = 0;
        memory[ 8284] = 1;
        memory[ 8285] = 0;
        memory[ 8286] = 0;
        memory[ 8287] = 0;
        memory[ 8288] = 1;
        memory[ 8289] = 0;
        memory[ 8290] = 1;
        memory[ 8291] = 0;
        memory[ 8292] = 0;
        memory[ 8293] = 0;
        memory[ 8294] = 0;
        memory[ 8295] = 0;
        memory[ 8296] = 0;
        memory[ 8297] = 0;
        memory[ 8298] = 0;
        memory[ 8299] = 0;
        memory[ 8300] = 0;
        memory[ 8301] = 1;
        memory[ 8302] = 0;
        memory[ 8303] = 0;
        memory[ 8304] = 0;
        memory[ 8305] = 0;
        memory[ 8306] = 1;
        memory[ 8307] = 0;
        memory[ 8308] = 0;
        memory[ 8309] = 1;
        memory[ 8310] = 0;
        memory[ 8311] = 0;
        memory[ 8312] = 0;
        memory[ 8313] = 0;
        memory[ 8314] = 0;
        memory[ 8315] = 0;
        memory[ 8316] = 0;
        memory[ 8317] = 0;
        memory[ 8318] = 0;
        memory[ 8319] = 0;
        memory[ 8320] = 0;
        memory[ 8321] = 0;
        memory[ 8322] = 0;
        memory[ 8323] = 0;
        memory[ 8324] = 1;
        memory[ 8325] = 0;
        memory[ 8326] = 0;
        memory[ 8327] = 1;
        memory[ 8328] = 1;
        memory[ 8329] = 0;
        memory[ 8330] = 0;
        memory[ 8331] = 1;
        memory[ 8332] = 0;
        memory[ 8333] = 0;
        memory[ 8334] = 0;
        memory[ 8335] = 0;
        memory[ 8336] = 0;
        memory[ 8337] = 0;
        memory[ 8338] = 0;
        memory[ 8339] = 0;
        memory[ 8340] = 0;
        memory[ 8341] = 0;
        memory[ 8342] = 0;
        memory[ 8343] = 0;
        memory[ 8344] = 0;
        memory[ 8345] = 0;
        memory[ 8346] = 1;
        memory[ 8347] = 1;
        memory[ 8348] = 0;
        memory[ 8349] = 0;
        memory[ 8350] = 0;
        memory[ 8351] = 0;
        memory[ 8352] = 0;
        memory[ 8353] = 0;
        memory[ 8354] = 0;
        memory[ 8355] = 0;
        memory[ 8356] = 0;
        memory[ 8357] = 0;
        memory[ 8358] = 0;
        memory[ 8359] = 0;
        memory[ 8360] = 1;
        memory[ 8361] = 0;
        memory[ 8362] = 1;
        memory[ 8363] = 0;
        memory[ 8364] = 0;
        memory[ 8365] = 0;
        memory[ 8366] = 0;
        memory[ 8367] = 0;
        memory[ 8368] = 0;
        memory[ 8369] = 0;
        memory[ 8370] = 0;
        memory[ 8371] = 0;
        memory[ 8372] = 0;
        memory[ 8373] = 0;
        memory[ 8374] = 0;
        memory[ 8375] = 0;
        memory[ 8376] = 1;
        memory[ 8377] = 0;
        memory[ 8378] = 0;
        memory[ 8379] = 0;
        memory[ 8380] = 0;
        memory[ 8381] = 0;
        memory[ 8382] = 0;
        memory[ 8383] = 0;
        memory[ 8384] = 0;
        memory[ 8385] = 0;
        memory[ 8386] = 0;
        memory[ 8387] = 0;
        memory[ 8388] = 0;
        memory[ 8389] = 0;
        memory[ 8390] = 0;
        memory[ 8391] = 0;
        memory[ 8392] = 0;
        memory[ 8393] = 1;
        memory[ 8394] = 0;
        memory[ 8395] = 0;
        memory[ 8396] = 1;
        memory[ 8397] = 1;
        memory[ 8398] = 0;
        memory[ 8399] = 0;
        memory[ 8400] = 0;
        memory[ 8401] = 0;
        memory[ 8402] = 0;
        memory[ 8403] = 0;
        memory[ 8404] = 1;
        memory[ 8405] = 0;
        memory[ 8406] = 0;
        memory[ 8407] = 0;
        memory[ 8408] = 0;
        memory[ 8409] = 0;
        memory[ 8410] = 0;
        memory[ 8411] = 0;
        memory[ 8412] = 0;
        memory[ 8413] = 0;
        memory[ 8414] = 0;
        memory[ 8415] = 0;
        memory[ 8416] = 0;
        memory[ 8417] = 0;
        memory[ 8418] = 1;
        memory[ 8419] = 0;
        memory[ 8420] = 1;
        memory[ 8421] = 1;
        memory[ 8422] = 1;
        memory[ 8423] = 0;
        memory[ 8424] = 1;
        memory[ 8425] = 0;
        memory[ 8426] = 0;
        memory[ 8427] = 0;
        memory[ 8428] = 0;
        memory[ 8429] = 0;
        memory[ 8430] = 0;
        memory[ 8431] = 0;
        memory[ 8432] = 0;
        memory[ 8433] = 0;
        memory[ 8434] = 0;
        memory[ 8435] = 0;
        memory[ 8436] = 0;
        memory[ 8437] = 0;
        memory[ 8438] = 1;
        memory[ 8439] = 0;
        memory[ 8440] = 0;
        memory[ 8441] = 0;
        memory[ 8442] = 0;
        memory[ 8443] = 0;
        memory[ 8444] = 0;
        memory[ 8445] = 0;
        memory[ 8446] = 0;
        memory[ 8447] = 0;
        memory[ 8448] = 0;
        memory[ 8449] = 0;
        memory[ 8450] = 0;
        memory[ 8451] = 0;
        memory[ 8452] = 0;
        memory[ 8453] = 1;
        memory[ 8454] = 1;
        memory[ 8455] = 1;
        memory[ 8456] = 0;
        memory[ 8457] = 0;
        memory[ 8458] = 0;
        memory[ 8459] = 0;
        memory[ 8460] = 0;
        memory[ 8461] = 0;
        memory[ 8462] = 0;
        memory[ 8463] = 0;
        memory[ 8464] = 0;
        memory[ 8465] = 0;
        memory[ 8466] = 0;
        memory[ 8467] = 0;
        memory[ 8468] = 0;
        memory[ 8469] = 0;
        memory[ 8470] = 0;
        memory[ 8471] = 0;
        memory[ 8472] = 0;
        memory[ 8473] = 0;
        memory[ 8474] = 0;
        memory[ 8475] = 0;
        memory[ 8476] = 1;
        memory[ 8477] = 0;
        memory[ 8478] = 0;
        memory[ 8479] = 0;
        memory[ 8480] = 0;
        memory[ 8481] = 1;
        memory[ 8482] = 0;
        memory[ 8483] = 0;
        memory[ 8484] = 0;
        memory[ 8485] = 0;
        memory[ 8486] = 0;
        memory[ 8487] = 1;
        memory[ 8488] = 1;
        memory[ 8489] = 0;
        memory[ 8490] = 0;
        memory[ 8491] = 0;
        memory[ 8492] = 0;
        memory[ 8493] = 0;
        memory[ 8494] = 0;
        memory[ 8495] = 0;
        memory[ 8496] = 0;
        memory[ 8497] = 0;
        memory[ 8498] = 0;
        memory[ 8499] = 0;
        memory[ 8500] = 0;
        memory[ 8501] = 0;
        memory[ 8502] = 0;
        memory[ 8503] = 1;
        memory[ 8504] = 0;
        memory[ 8505] = 1;
        memory[ 8506] = 1;
        memory[ 8507] = 0;
        memory[ 8508] = 0;
        memory[ 8509] = 0;
        memory[ 8510] = 0;
        memory[ 8511] = 0;
        memory[ 8512] = 0;
        memory[ 8513] = 0;
        memory[ 8514] = 0;
        memory[ 8515] = 0;
        memory[ 8516] = 0;
        memory[ 8517] = 0;
        memory[ 8518] = 0;
        memory[ 8519] = 0;
        memory[ 8520] = 0;
        memory[ 8521] = 0;
        memory[ 8522] = 0;
        memory[ 8523] = 0;
        memory[ 8524] = 1;
        memory[ 8525] = 1;
        memory[ 8526] = 0;
        memory[ 8527] = 1;
        memory[ 8528] = 1;
        memory[ 8529] = 0;
        memory[ 8530] = 1;
        memory[ 8531] = 1;
        memory[ 8532] = 0;
        memory[ 8533] = 0;
        memory[ 8534] = 0;
        memory[ 8535] = 0;
        memory[ 8536] = 0;
        memory[ 8537] = 0;
        memory[ 8538] = 0;
        memory[ 8539] = 0;
        memory[ 8540] = 0;
        memory[ 8541] = 0;
        memory[ 8542] = 0;
        memory[ 8543] = 0;
        memory[ 8544] = 0;
        memory[ 8545] = 0;
        memory[ 8546] = 0;
        memory[ 8547] = 0;
        memory[ 8548] = 0;
        memory[ 8549] = 1;
        memory[ 8550] = 0;
        memory[ 8551] = 0;
        memory[ 8552] = 0;
        memory[ 8553] = 0;
        memory[ 8554] = 0;
        memory[ 8555] = 0;
        memory[ 8556] = 0;
        memory[ 8557] = 0;
        memory[ 8558] = 1;
        memory[ 8559] = 0;
        memory[ 8560] = 0;
        memory[ 8561] = 0;
        memory[ 8562] = 0;
        memory[ 8563] = 0;
        memory[ 8564] = 0;
        memory[ 8565] = 0;
        memory[ 8566] = 0;
        memory[ 8567] = 1;
        memory[ 8568] = 1;
        memory[ 8569] = 0;
        memory[ 8570] = 0;
        memory[ 8571] = 1;
        memory[ 8572] = 0;
        memory[ 8573] = 0;
        memory[ 8574] = 0;
        memory[ 8575] = 0;
        memory[ 8576] = 0;
        memory[ 8577] = 0;
        memory[ 8578] = 0;
        memory[ 8579] = 0;
        memory[ 8580] = 0;
        memory[ 8581] = 0;
        memory[ 8582] = 0;
        memory[ 8583] = 1;
        memory[ 8584] = 1;
        memory[ 8585] = 0;
        memory[ 8586] = 0;
        memory[ 8587] = 0;
        memory[ 8588] = 0;
        memory[ 8589] = 0;
        memory[ 8590] = 1;
        memory[ 8591] = 1;
        memory[ 8592] = 1;
        memory[ 8593] = 0;
        memory[ 8594] = 1;
        memory[ 8595] = 0;
        memory[ 8596] = 0;
        memory[ 8597] = 0;
        memory[ 8598] = 0;
        memory[ 8599] = 0;
        memory[ 8600] = 0;
        memory[ 8601] = 0;
        memory[ 8602] = 0;
        memory[ 8603] = 0;
        memory[ 8604] = 0;
        memory[ 8605] = 0;
        memory[ 8606] = 0;
        memory[ 8607] = 0;
        memory[ 8608] = 0;
        memory[ 8609] = 0;
        memory[ 8610] = 0;
        memory[ 8611] = 0;
        memory[ 8612] = 0;
        memory[ 8613] = 0;
        memory[ 8614] = 0;
        memory[ 8615] = 0;
        memory[ 8616] = 1;
        memory[ 8617] = 0;
        memory[ 8618] = 1;
        memory[ 8619] = 0;
        memory[ 8620] = 1;
        memory[ 8621] = 0;
        memory[ 8622] = 0;
        memory[ 8623] = 0;
        memory[ 8624] = 0;
        memory[ 8625] = 1;
        memory[ 8626] = 0;
        memory[ 8627] = 0;
        memory[ 8628] = 0;
        memory[ 8629] = 0;
        memory[ 8630] = 0;
        memory[ 8631] = 0;
        memory[ 8632] = 0;
        memory[ 8633] = 0;
        memory[ 8634] = 0;
        memory[ 8635] = 0;
        memory[ 8636] = 0;
        memory[ 8637] = 0;
        memory[ 8638] = 0;
        memory[ 8639] = 0;
        memory[ 8640] = 0;
        memory[ 8641] = 0;
        memory[ 8642] = 0;
        memory[ 8643] = 0;
        memory[ 8644] = 0;
        memory[ 8645] = 0;
        memory[ 8646] = 0;
        memory[ 8647] = 0;
        memory[ 8648] = 0;
        memory[ 8649] = 0;
        memory[ 8650] = 0;
        memory[ 8651] = 0;
        memory[ 8652] = 0;
        memory[ 8653] = 0;
        memory[ 8654] = 0;
        memory[ 8655] = 1;
        memory[ 8656] = 0;
        memory[ 8657] = 0;
        memory[ 8658] = 0;
        memory[ 8659] = 1;
        memory[ 8660] = 0;
        memory[ 8661] = 0;
        memory[ 8662] = 0;
        memory[ 8663] = 0;
        memory[ 8664] = 0;
        memory[ 8665] = 0;
        memory[ 8666] = 0;
        memory[ 8667] = 0;
        memory[ 8668] = 0;
        memory[ 8669] = 0;
        memory[ 8670] = 0;
        memory[ 8671] = 0;
        memory[ 8672] = 0;
        memory[ 8673] = 0;
        memory[ 8674] = 1;
        memory[ 8675] = 1;
        memory[ 8676] = 0;
        memory[ 8677] = 0;
        memory[ 8678] = 0;
        memory[ 8679] = 0;
        memory[ 8680] = 0;
        memory[ 8681] = 0;
        memory[ 8682] = 1;
        memory[ 8683] = 0;
        memory[ 8684] = 0;
        memory[ 8685] = 0;
        memory[ 8686] = 0;
        memory[ 8687] = 0;
        memory[ 8688] = 0;
        memory[ 8689] = 0;
        memory[ 8690] = 0;
        memory[ 8691] = 0;
        memory[ 8692] = 0;
        memory[ 8693] = 0;
        memory[ 8694] = 0;
        memory[ 8695] = 0;
        memory[ 8696] = 1;
        memory[ 8697] = 1;
        memory[ 8698] = 1;
        memory[ 8699] = 1;
        memory[ 8700] = 0;
        memory[ 8701] = 0;
        memory[ 8702] = 0;
        memory[ 8703] = 0;
        memory[ 8704] = 0;
        memory[ 8705] = 1;
        memory[ 8706] = 0;
        memory[ 8707] = 0;
        memory[ 8708] = 0;
        memory[ 8709] = 0;
        memory[ 8710] = 0;
        memory[ 8711] = 0;
        memory[ 8712] = 0;
        memory[ 8713] = 0;
        memory[ 8714] = 1;
        memory[ 8715] = 1;
        memory[ 8716] = 0;
        memory[ 8717] = 0;
        memory[ 8718] = 0;
        memory[ 8719] = 1;
        memory[ 8720] = 1;
        memory[ 8721] = 0;
        memory[ 8722] = 0;
        memory[ 8723] = 0;
        memory[ 8724] = 0;
        memory[ 8725] = 0;
        memory[ 8726] = 0;
        memory[ 8727] = 0;
        memory[ 8728] = 1;
        memory[ 8729] = 1;
        memory[ 8730] = 1;
        memory[ 8731] = 0;
        memory[ 8732] = 0;
        memory[ 8733] = 0;
        memory[ 8734] = 0;
        memory[ 8735] = 0;
        memory[ 8736] = 0;
        memory[ 8737] = 0;
        memory[ 8738] = 0;
        memory[ 8739] = 0;
        memory[ 8740] = 0;
        memory[ 8741] = 0;
        memory[ 8742] = 0;
        memory[ 8743] = 0;
        memory[ 8744] = 0;
        memory[ 8745] = 0;
        memory[ 8746] = 0;
        memory[ 8747] = 0;
        memory[ 8748] = 0;
        memory[ 8749] = 0;
        memory[ 8750] = 0;
        memory[ 8751] = 0;
        memory[ 8752] = 0;
        memory[ 8753] = 0;
        memory[ 8754] = 0;
        memory[ 8755] = 0;
        memory[ 8756] = 0;
        memory[ 8757] = 0;
        memory[ 8758] = 0;
        memory[ 8759] = 0;
        memory[ 8760] = 0;
        memory[ 8761] = 0;
        memory[ 8762] = 1;
        memory[ 8763] = 1;
        memory[ 8764] = 1;
        memory[ 8765] = 0;
        memory[ 8766] = 1;
        memory[ 8767] = 0;
        memory[ 8768] = 0;
        memory[ 8769] = 1;
        memory[ 8770] = 1;
        memory[ 8771] = 1;
        memory[ 8772] = 0;
        memory[ 8773] = 0;
        memory[ 8774] = 0;
        memory[ 8775] = 0;
        memory[ 8776] = 0;
        memory[ 8777] = 0;
        memory[ 8778] = 0;
        memory[ 8779] = 0;
        memory[ 8780] = 0;
        memory[ 8781] = 1;
        memory[ 8782] = 1;
        memory[ 8783] = 0;
        memory[ 8784] = 0;
        memory[ 8785] = 0;
        memory[ 8786] = 0;
        memory[ 8787] = 0;
        memory[ 8788] = 0;
        memory[ 8789] = 0;
        memory[ 8790] = 0;
        memory[ 8791] = 0;
        memory[ 8792] = 0;
        memory[ 8793] = 0;
        memory[ 8794] = 0;
        memory[ 8795] = 0;
        memory[ 8796] = 0;
        memory[ 8797] = 0;
        memory[ 8798] = 0;
        memory[ 8799] = 0;
        memory[ 8800] = 0;
        memory[ 8801] = 0;
        memory[ 8802] = 1;
        memory[ 8803] = 1;
        memory[ 8804] = 0;
        memory[ 8805] = 1;
        memory[ 8806] = 0;
        memory[ 8807] = 0;
        memory[ 8808] = 0;
        memory[ 8809] = 0;
        memory[ 8810] = 0;
        memory[ 8811] = 0;
        memory[ 8812] = 0;
        memory[ 8813] = 0;
        memory[ 8814] = 0;
        memory[ 8815] = 0;
        memory[ 8816] = 0;
        memory[ 8817] = 0;
        memory[ 8818] = 0;
        memory[ 8819] = 0;
        memory[ 8820] = 0;
        memory[ 8821] = 0;
        memory[ 8822] = 0;
        memory[ 8823] = 0;
        memory[ 8824] = 0;
        memory[ 8825] = 0;
        memory[ 8826] = 0;
        memory[ 8827] = 0;
        memory[ 8828] = 0;
        memory[ 8829] = 0;
        memory[ 8830] = 0;
        memory[ 8831] = 0;
        memory[ 8832] = 0;
        memory[ 8833] = 0;
        memory[ 8834] = 0;
        memory[ 8835] = 0;
        memory[ 8836] = 0;
        memory[ 8837] = 0;
        memory[ 8838] = 0;
        memory[ 8839] = 0;
        memory[ 8840] = 0;
        memory[ 8841] = 0;
        memory[ 8842] = 0;
        memory[ 8843] = 0;
        memory[ 8844] = 1;
        memory[ 8845] = 0;
        memory[ 8846] = 0;
        memory[ 8847] = 0;
        memory[ 8848] = 0;
        memory[ 8849] = 1;
        memory[ 8850] = 0;
        memory[ 8851] = 0;
        memory[ 8852] = 0;
        memory[ 8853] = 0;
        memory[ 8854] = 0;
        memory[ 8855] = 0;
        memory[ 8856] = 0;
        memory[ 8857] = 0;
        memory[ 8858] = 0;
        memory[ 8859] = 0;
        memory[ 8860] = 0;
        memory[ 8861] = 0;
        memory[ 8862] = 0;
        memory[ 8863] = 0;
        memory[ 8864] = 0;
        memory[ 8865] = 0;
        memory[ 8866] = 0;
        memory[ 8867] = 0;
        memory[ 8868] = 0;
        memory[ 8869] = 0;
        memory[ 8870] = 0;
        memory[ 8871] = 0;
        memory[ 8872] = 0;
        memory[ 8873] = 0;
        memory[ 8874] = 0;
        memory[ 8875] = 0;
        memory[ 8876] = 0;
        memory[ 8877] = 0;
        memory[ 8878] = 0;
        memory[ 8879] = 0;
        memory[ 8880] = 1;
        memory[ 8881] = 0;
        memory[ 8882] = 0;
        memory[ 8883] = 0;
        memory[ 8884] = 0;
        memory[ 8885] = 0;
        memory[ 8886] = 0;
        memory[ 8887] = 0;
        memory[ 8888] = 0;
        memory[ 8889] = 0;
        memory[ 8890] = 0;
        memory[ 8891] = 0;
        memory[ 8892] = 0;
        memory[ 8893] = 0;
        memory[ 8894] = 0;
        memory[ 8895] = 1;
        memory[ 8896] = 0;
        memory[ 8897] = 1;
        memory[ 8898] = 0;
        memory[ 8899] = 0;
        memory[ 8900] = 0;
        memory[ 8901] = 0;
        memory[ 8902] = 0;
        memory[ 8903] = 1;
        memory[ 8904] = 0;
        memory[ 8905] = 0;
        memory[ 8906] = 0;
        memory[ 8907] = 0;
        memory[ 8908] = 0;
        memory[ 8909] = 0;
        memory[ 8910] = 0;
        memory[ 8911] = 0;
        memory[ 8912] = 0;
        memory[ 8913] = 0;
        memory[ 8914] = 0;
        memory[ 8915] = 0;
        memory[ 8916] = 0;
        memory[ 8917] = 0;
        memory[ 8918] = 0;
        memory[ 8919] = 0;
        memory[ 8920] = 0;
        memory[ 8921] = 0;
        memory[ 8922] = 0;
        memory[ 8923] = 0;
        memory[ 8924] = 0;
        memory[ 8925] = 0;
        memory[ 8926] = 0;
        memory[ 8927] = 0;
        memory[ 8928] = 0;
        memory[ 8929] = 1;
        memory[ 8930] = 1;
        memory[ 8931] = 0;
        memory[ 8932] = 0;
        memory[ 8933] = 0;
        memory[ 8934] = 1;
        memory[ 8935] = 0;
        memory[ 8936] = 0;
        memory[ 8937] = 1;
        memory[ 8938] = 0;
        memory[ 8939] = 0;
        memory[ 8940] = 0;
        memory[ 8941] = 0;
        memory[ 8942] = 0;
        memory[ 8943] = 0;
        memory[ 8944] = 0;
        memory[ 8945] = 0;
        memory[ 8946] = 0;
        memory[ 8947] = 0;
        memory[ 8948] = 0;
        memory[ 8949] = 0;
        memory[ 8950] = 0;
        memory[ 8951] = 0;
        memory[ 8952] = 1;
        memory[ 8953] = 0;
        memory[ 8954] = 0;
        memory[ 8955] = 0;
        memory[ 8956] = 1;
        memory[ 8957] = 0;
        memory[ 8958] = 0;
        memory[ 8959] = 0;
        memory[ 8960] = 0;
        memory[ 8961] = 0;
        memory[ 8962] = 0;
        memory[ 8963] = 1;
        memory[ 8964] = 0;
        memory[ 8965] = 0;
        memory[ 8966] = 0;
        memory[ 8967] = 0;
        memory[ 8968] = 0;
        memory[ 8969] = 0;
        memory[ 8970] = 0;
        memory[ 8971] = 0;
        memory[ 8972] = 0;
        memory[ 8973] = 0;
        memory[ 8974] = 0;
        memory[ 8975] = 0;
        memory[ 8976] = 0;
        memory[ 8977] = 0;
        memory[ 8978] = 0;
        memory[ 8979] = 0;
        memory[ 8980] = 0;
        memory[ 8981] = 0;
        memory[ 8982] = 0;
        memory[ 8983] = 0;
        memory[ 8984] = 0;
        memory[ 8985] = 0;
        memory[ 8986] = 0;
        memory[ 8987] = 0;
        memory[ 8988] = 1;
        memory[ 8989] = 1;
        memory[ 8990] = 0;
        memory[ 8991] = 0;
        memory[ 8992] = 0;
        memory[ 8993] = 0;
        memory[ 8994] = 0;
        memory[ 8995] = 0;
        memory[ 8996] = 0;
        memory[ 8997] = 0;
        memory[ 8998] = 0;
        memory[ 8999] = 1;
        memory[ 9000] = 0;
        memory[ 9001] = 0;
        memory[ 9002] = 1;
        memory[ 9003] = 0;
        memory[ 9004] = 0;
        memory[ 9005] = 0;
        memory[ 9006] = 0;
        memory[ 9007] = 0;
        memory[ 9008] = 0;
        memory[ 9009] = 0;
        memory[ 9010] = 0;
        memory[ 9011] = 0;
        memory[ 9012] = 0;
        memory[ 9013] = 0;
        memory[ 9014] = 0;
        memory[ 9015] = 0;
        memory[ 9016] = 0;
        memory[ 9017] = 0;
        memory[ 9018] = 0;
        memory[ 9019] = 0;
        memory[ 9020] = 0;
        memory[ 9021] = 0;
        memory[ 9022] = 0;
        memory[ 9023] = 1;
        memory[ 9024] = 0;
        memory[ 9025] = 0;
        memory[ 9026] = 0;
        memory[ 9027] = 0;
        memory[ 9028] = 0;
        memory[ 9029] = 0;
        memory[ 9030] = 0;
        memory[ 9031] = 0;
        memory[ 9032] = 0;
        memory[ 9033] = 0;
        memory[ 9034] = 0;
        memory[ 9035] = 0;
        memory[ 9036] = 0;
        memory[ 9037] = 0;
        memory[ 9038] = 0;
        memory[ 9039] = 0;
        memory[ 9040] = 0;
        memory[ 9041] = 0;
        memory[ 9042] = 0;
        memory[ 9043] = 0;
        memory[ 9044] = 0;
        memory[ 9045] = 0;
        memory[ 9046] = 0;
        memory[ 9047] = 0;
        memory[ 9048] = 0;
        memory[ 9049] = 0;
        memory[ 9050] = 0;
        memory[ 9051] = 0;
        memory[ 9052] = 0;
        memory[ 9053] = 0;
        memory[ 9054] = 0;
        memory[ 9055] = 0;
        memory[ 9056] = 0;
        memory[ 9057] = 0;
        memory[ 9058] = 0;
        memory[ 9059] = 0;
        memory[ 9060] = 0;
        memory[ 9061] = 0;
        memory[ 9062] = 0;
        memory[ 9063] = 0;
        memory[ 9064] = 0;
        memory[ 9065] = 0;
        memory[ 9066] = 0;
        memory[ 9067] = 0;
        memory[ 9068] = 0;
        memory[ 9069] = 0;
        memory[ 9070] = 0;
        memory[ 9071] = 0;
        memory[ 9072] = 0;
        memory[ 9073] = 0;
        memory[ 9074] = 0;
        memory[ 9075] = 1;
        memory[ 9076] = 0;
        memory[ 9077] = 0;
        memory[ 9078] = 0;
        memory[ 9079] = 0;
        memory[ 9080] = 1;
        memory[ 9081] = 0;
        memory[ 9082] = 0;
        memory[ 9083] = 1;
        memory[ 9084] = 0;
        memory[ 9085] = 0;
        memory[ 9086] = 0;
        memory[ 9087] = 0;
        memory[ 9088] = 0;
        memory[ 9089] = 0;
        memory[ 9090] = 0;
        memory[ 9091] = 0;
        memory[ 9092] = 0;
        memory[ 9093] = 0;
        memory[ 9094] = 0;
        memory[ 9095] = 0;
        memory[ 9096] = 0;
        memory[ 9097] = 0;
        memory[ 9098] = 0;
        memory[ 9099] = 0;
        memory[ 9100] = 0;
        memory[ 9101] = 0;
        memory[ 9102] = 0;
        memory[ 9103] = 0;
        memory[ 9104] = 0;
        memory[ 9105] = 0;
        memory[ 9106] = 0;
        memory[ 9107] = 0;
        memory[ 9108] = 0;
        memory[ 9109] = 0;
        memory[ 9110] = 0;
        memory[ 9111] = 0;
        memory[ 9112] = 0;
        memory[ 9113] = 1;
        memory[ 9114] = 0;
        memory[ 9115] = 0;
        memory[ 9116] = 0;
        memory[ 9117] = 0;
        memory[ 9118] = 0;
        memory[ 9119] = 0;
        memory[ 9120] = 0;
        memory[ 9121] = 0;
        memory[ 9122] = 0;
        memory[ 9123] = 0;
        memory[ 9124] = 0;
        memory[ 9125] = 0;
        memory[ 9126] = 0;
        memory[ 9127] = 0;
        memory[ 9128] = 0;
        memory[ 9129] = 0;
        memory[ 9130] = 1;
        memory[ 9131] = 0;
        memory[ 9132] = 0;
        memory[ 9133] = 0;
        memory[ 9134] = 0;
        memory[ 9135] = 0;
        memory[ 9136] = 0;
        memory[ 9137] = 0;
        memory[ 9138] = 0;
        memory[ 9139] = 0;
        memory[ 9140] = 0;
        memory[ 9141] = 0;
        memory[ 9142] = 0;
        memory[ 9143] = 0;
        memory[ 9144] = 0;
        memory[ 9145] = 0;
        memory[ 9146] = 1;
        memory[ 9147] = 0;
        memory[ 9148] = 0;
        memory[ 9149] = 0;
        memory[ 9150] = 0;
        memory[ 9151] = 0;
        memory[ 9152] = 0;
        memory[ 9153] = 0;
        memory[ 9154] = 0;
        memory[ 9155] = 0;
        memory[ 9156] = 0;
        memory[ 9157] = 0;
        memory[ 9158] = 0;
        memory[ 9159] = 0;
        memory[ 9160] = 0;
        memory[ 9161] = 0;
        memory[ 9162] = 0;
        memory[ 9163] = 0;
        memory[ 9164] = 0;
        memory[ 9165] = 0;
        memory[ 9166] = 0;
        memory[ 9167] = 0;
        memory[ 9168] = 0;
        memory[ 9169] = 0;
        memory[ 9170] = 0;
        memory[ 9171] = 0;
        memory[ 9172] = 0;
        memory[ 9173] = 0;
        memory[ 9174] = 0;
        memory[ 9175] = 0;
        memory[ 9176] = 0;
        memory[ 9177] = 0;
        memory[ 9178] = 0;
        memory[ 9179] = 0;
        memory[ 9180] = 0;
        memory[ 9181] = 0;
        memory[ 9182] = 0;
        memory[ 9183] = 0;
        memory[ 9184] = 0;
        memory[ 9185] = 0;
        memory[ 9186] = 0;
        memory[ 9187] = 0;
        memory[ 9188] = 0;
        memory[ 9189] = 0;
        memory[ 9190] = 0;
        memory[ 9191] = 0;
        memory[ 9192] = 1;
        memory[ 9193] = 0;
        memory[ 9194] = 0;
        memory[ 9195] = 0;
        memory[ 9196] = 1;
        memory[ 9197] = 0;
        memory[ 9198] = 0;
        memory[ 9199] = 0;
        memory[ 9200] = 0;
        memory[ 9201] = 0;
        memory[ 9202] = 0;
        memory[ 9203] = 0;
        memory[ 9204] = 0;
        memory[ 9205] = 0;
        memory[ 9206] = 0;
        memory[ 9207] = 0;
        memory[ 9208] = 1;
        memory[ 9209] = 0;
        memory[ 9210] = 0;
        memory[ 9211] = 1;
        memory[ 9212] = 0;
        memory[ 9213] = 0;
        memory[ 9214] = 0;
        memory[ 9215] = 0;
        memory[ 9216] = 0;
        memory[ 9217] = 0;
        memory[ 9218] = 0;
        memory[ 9219] = 0;
        memory[ 9220] = 0;
        memory[ 9221] = 0;
        memory[ 9222] = 0;
        memory[ 9223] = 0;
        memory[ 9224] = 0;
        memory[ 9225] = 0;
        memory[ 9226] = 0;
        memory[ 9227] = 0;
        memory[ 9228] = 0;
        memory[ 9229] = 0;
        memory[ 9230] = 0;
        memory[ 9231] = 0;
        memory[ 9232] = 0;
        memory[ 9233] = 0;
        memory[ 9234] = 0;
        memory[ 9235] = 0;
        memory[ 9236] = 0;
        memory[ 9237] = 0;
        memory[ 9238] = 0;
        memory[ 9239] = 0;
        memory[ 9240] = 0;
        memory[ 9241] = 0;
        memory[ 9242] = 0;
        memory[ 9243] = 0;
        memory[ 9244] = 0;
        memory[ 9245] = 0;
        memory[ 9246] = 0;
        memory[ 9247] = 0;
        memory[ 9248] = 0;
        memory[ 9249] = 0;
        memory[ 9250] = 0;
        memory[ 9251] = 0;
        memory[ 9252] = 0;
        memory[ 9253] = 0;
        memory[ 9254] = 0;
        memory[ 9255] = 0;
        memory[ 9256] = 0;
        memory[ 9257] = 0;
        memory[ 9258] = 0;
        memory[ 9259] = 0;
        memory[ 9260] = 0;
        memory[ 9261] = 0;
        memory[ 9262] = 0;
        memory[ 9263] = 0;
        memory[ 9264] = 0;
        memory[ 9265] = 0;
        memory[ 9266] = 0;
        memory[ 9267] = 0;
        memory[ 9268] = 0;
        memory[ 9269] = 0;
        memory[ 9270] = 0;
        memory[ 9271] = 0;
        memory[ 9272] = 0;
        memory[ 9273] = 0;
        memory[ 9274] = 0;
        memory[ 9275] = 0;
        memory[ 9276] = 0;
        memory[ 9277] = 1;
        memory[ 9278] = 0;
        memory[ 9279] = 0;
        memory[ 9280] = 0;
        memory[ 9281] = 0;
        memory[ 9282] = 0;
        memory[ 9283] = 1;
        memory[ 9284] = 0;
        memory[ 9285] = 0;
        memory[ 9286] = 0;
        memory[ 9287] = 0;
        memory[ 9288] = 0;
        memory[ 9289] = 0;
        memory[ 9290] = 0;
        memory[ 9291] = 0;
        memory[ 9292] = 0;
        memory[ 9293] = 1;
        memory[ 9294] = 0;
        memory[ 9295] = 0;
        memory[ 9296] = 0;
        memory[ 9297] = 1;
        memory[ 9298] = 0;
        memory[ 9299] = 0;
        memory[ 9300] = 0;
        memory[ 9301] = 0;
        memory[ 9302] = 0;
        memory[ 9303] = 0;
        memory[ 9304] = 0;
        memory[ 9305] = 0;
        memory[ 9306] = 0;
        memory[ 9307] = 0;
        memory[ 9308] = 1;
        memory[ 9309] = 1;
        memory[ 9310] = 0;
        memory[ 9311] = 1;
        memory[ 9312] = 0;
        memory[ 9313] = 0;
        memory[ 9314] = 1;
        memory[ 9315] = 0;
        memory[ 9316] = 0;
        memory[ 9317] = 1;
        memory[ 9318] = 1;
        memory[ 9319] = 0;
        memory[ 9320] = 0;
        memory[ 9321] = 0;
        memory[ 9322] = 0;
        memory[ 9323] = 0;
        memory[ 9324] = 0;
        memory[ 9325] = 0;
        memory[ 9326] = 0;
        memory[ 9327] = 0;
        memory[ 9328] = 0;
        memory[ 9329] = 0;
        memory[ 9330] = 0;
        memory[ 9331] = 0;
        memory[ 9332] = 0;
        memory[ 9333] = 0;
        memory[ 9334] = 0;
        memory[ 9335] = 0;
        memory[ 9336] = 0;
        memory[ 9337] = 0;
        memory[ 9338] = 0;
        memory[ 9339] = 0;
        memory[ 9340] = 0;
        memory[ 9341] = 0;
        memory[ 9342] = 0;
        memory[ 9343] = 0;
        memory[ 9344] = 0;
        memory[ 9345] = 0;
        memory[ 9346] = 0;
        memory[ 9347] = 1;
        memory[ 9348] = 0;
        memory[ 9349] = 0;
        memory[ 9350] = 0;
        memory[ 9351] = 0;
        memory[ 9352] = 0;
        memory[ 9353] = 0;
        memory[ 9354] = 0;
        memory[ 9355] = 0;
        memory[ 9356] = 0;
        memory[ 9357] = 0;
        memory[ 9358] = 0;
        memory[ 9359] = 0;
        memory[ 9360] = 0;
        memory[ 9361] = 0;
        memory[ 9362] = 0;
        memory[ 9363] = 0;
        memory[ 9364] = 0;
        memory[ 9365] = 0;
        memory[ 9366] = 1;
        memory[ 9367] = 1;
        memory[ 9368] = 0;
        memory[ 9369] = 0;
        memory[ 9370] = 0;
        memory[ 9371] = 0;
        memory[ 9372] = 0;
        memory[ 9373] = 0;
        memory[ 9374] = 0;
        memory[ 9375] = 0;
        memory[ 9376] = 0;
        memory[ 9377] = 0;
        memory[ 9378] = 0;
        memory[ 9379] = 0;
        memory[ 9380] = 0;
        memory[ 9381] = 0;
        memory[ 9382] = 0;
        memory[ 9383] = 0;
        memory[ 9384] = 0;
        memory[ 9385] = 0;
        memory[ 9386] = 0;
        memory[ 9387] = 0;
        memory[ 9388] = 0;
        memory[ 9389] = 0;
        memory[ 9390] = 1;
        memory[ 9391] = 0;
        memory[ 9392] = 0;
        memory[ 9393] = 0;
        memory[ 9394] = 0;
        memory[ 9395] = 0;
        memory[ 9396] = 0;
        memory[ 9397] = 0;
        memory[ 9398] = 0;
        memory[ 9399] = 0;
        memory[ 9400] = 1;
        memory[ 9401] = 0;
        memory[ 9402] = 0;
        memory[ 9403] = 0;
        memory[ 9404] = 0;
        memory[ 9405] = 0;
        memory[ 9406] = 0;
        memory[ 9407] = 0;
        memory[ 9408] = 0;
        memory[ 9409] = 0;
        memory[ 9410] = 0;
        memory[ 9411] = 0;
        memory[ 9412] = 1;
        memory[ 9413] = 1;
        memory[ 9414] = 1;
        memory[ 9415] = 1;
        memory[ 9416] = 0;
        memory[ 9417] = 0;
        memory[ 9418] = 0;
        memory[ 9419] = 0;
        memory[ 9420] = 1;
        memory[ 9421] = 0;
        memory[ 9422] = 0;
        memory[ 9423] = 0;
        memory[ 9424] = 0;
        memory[ 9425] = 1;
        memory[ 9426] = 0;
        memory[ 9427] = 0;
        memory[ 9428] = 0;
        memory[ 9429] = 0;
        memory[ 9430] = 0;
        memory[ 9431] = 0;
        memory[ 9432] = 0;
        memory[ 9433] = 0;
        memory[ 9434] = 0;
        memory[ 9435] = 0;
        memory[ 9436] = 0;
        memory[ 9437] = 0;
        memory[ 9438] = 0;
        memory[ 9439] = 0;
        memory[ 9440] = 0;
        memory[ 9441] = 0;
        memory[ 9442] = 0;
        memory[ 9443] = 1;
        memory[ 9444] = 0;
        memory[ 9445] = 0;
        memory[ 9446] = 0;
        memory[ 9447] = 0;
        memory[ 9448] = 0;
        memory[ 9449] = 0;
        memory[ 9450] = 0;
        memory[ 9451] = 0;
        memory[ 9452] = 0;
        memory[ 9453] = 0;
        memory[ 9454] = 0;
        memory[ 9455] = 0;
        memory[ 9456] = 0;
        memory[ 9457] = 0;
        memory[ 9458] = 0;
        memory[ 9459] = 0;
        memory[ 9460] = 0;
        memory[ 9461] = 0;
        memory[ 9462] = 0;
        memory[ 9463] = 0;
        memory[ 9464] = 0;
        memory[ 9465] = 0;
        memory[ 9466] = 0;
        memory[ 9467] = 0;
        memory[ 9468] = 0;
        memory[ 9469] = 0;
        memory[ 9470] = 0;
        memory[ 9471] = 0;
        memory[ 9472] = 0;
        memory[ 9473] = 0;
        memory[ 9474] = 1;
        memory[ 9475] = 0;
        memory[ 9476] = 0;
        memory[ 9477] = 1;
        memory[ 9478] = 0;
        memory[ 9479] = 0;
        memory[ 9480] = 0;
        memory[ 9481] = 0;
        memory[ 9482] = 0;
        memory[ 9483] = 0;
        memory[ 9484] = 1;
        memory[ 9485] = 0;
        memory[ 9486] = 0;
        memory[ 9487] = 0;
        memory[ 9488] = 0;
        memory[ 9489] = 0;
        memory[ 9490] = 0;
        memory[ 9491] = 0;
        memory[ 9492] = 0;
        memory[ 9493] = 0;
        memory[ 9494] = 0;
        memory[ 9495] = 0;
        memory[ 9496] = 0;
        memory[ 9497] = 0;
        memory[ 9498] = 0;
        memory[ 9499] = 0;
        memory[ 9500] = 0;
        memory[ 9501] = 1;
        memory[ 9502] = 0;
        memory[ 9503] = 0;
        memory[ 9504] = 1;
        memory[ 9505] = 0;
        memory[ 9506] = 0;
        memory[ 9507] = 0;
        memory[ 9508] = 0;
        memory[ 9509] = 0;
        memory[ 9510] = 0;
        memory[ 9511] = 0;
        memory[ 9512] = 0;
        memory[ 9513] = 0;
        memory[ 9514] = 0;
        memory[ 9515] = 0;
        memory[ 9516] = 0;
        memory[ 9517] = 0;
        memory[ 9518] = 1;
        memory[ 9519] = 1;
        memory[ 9520] = 1;
        memory[ 9521] = 0;
        memory[ 9522] = 0;
        memory[ 9523] = 0;
        memory[ 9524] = 0;
        memory[ 9525] = 0;
        memory[ 9526] = 0;
        memory[ 9527] = 0;
        memory[ 9528] = 0;
        memory[ 9529] = 0;
        memory[ 9530] = 0;
        memory[ 9531] = 0;
        memory[ 9532] = 1;
        memory[ 9533] = 1;
        memory[ 9534] = 1;
        memory[ 9535] = 0;
        memory[ 9536] = 0;
        memory[ 9537] = 0;
        memory[ 9538] = 0;
        memory[ 9539] = 0;
        memory[ 9540] = 0;
        memory[ 9541] = 0;
        memory[ 9542] = 0;
        memory[ 9543] = 0;
        memory[ 9544] = 0;
        memory[ 9545] = 0;
        memory[ 9546] = 0;
        memory[ 9547] = 1;
        memory[ 9548] = 0;
        memory[ 9549] = 0;
        memory[ 9550] = 0;
        memory[ 9551] = 1;
        memory[ 9552] = 1;
        memory[ 9553] = 0;
        memory[ 9554] = 0;
        memory[ 9555] = 0;
        memory[ 9556] = 0;
        memory[ 9557] = 0;
        memory[ 9558] = 0;
        memory[ 9559] = 0;
        memory[ 9560] = 0;
        memory[ 9561] = 0;
        memory[ 9562] = 0;
        memory[ 9563] = 0;
        memory[ 9564] = 0;
        memory[ 9565] = 0;
        memory[ 9566] = 0;
        memory[ 9567] = 0;
        memory[ 9568] = 0;
        memory[ 9569] = 0;
        memory[ 9570] = 0;
        memory[ 9571] = 0;
        memory[ 9572] = 0;
        memory[ 9573] = 0;
        memory[ 9574] = 0;
        memory[ 9575] = 0;
        memory[ 9576] = 0;
        memory[ 9577] = 0;
        memory[ 9578] = 0;
        memory[ 9579] = 0;
        memory[ 9580] = 0;
        memory[ 9581] = 0;
        memory[ 9582] = 0;
        memory[ 9583] = 0;
        memory[ 9584] = 0;
        memory[ 9585] = 0;
        memory[ 9586] = 0;
        memory[ 9587] = 0;
        memory[ 9588] = 1;
        memory[ 9589] = 0;
        memory[ 9590] = 0;
        memory[ 9591] = 1;
        memory[ 9592] = 0;
        memory[ 9593] = 0;
        memory[ 9594] = 0;
        memory[ 9595] = 0;
        memory[ 9596] = 0;
        memory[ 9597] = 1;
        memory[ 9598] = 0;
        memory[ 9599] = 0;
        memory[ 9600] = 0;
        memory[ 9601] = 0;
        memory[ 9602] = 0;
        memory[ 9603] = 0;
        memory[ 9604] = 0;
        memory[ 9605] = 1;
        memory[ 9606] = 1;
        memory[ 9607] = 1;
        memory[ 9608] = 0;
        memory[ 9609] = 0;
        memory[ 9610] = 0;
        memory[ 9611] = 0;
        memory[ 9612] = 0;
        memory[ 9613] = 0;
        memory[ 9614] = 1;
        memory[ 9615] = 1;
        memory[ 9616] = 0;
        memory[ 9617] = 0;
        memory[ 9618] = 0;
        memory[ 9619] = 0;
        memory[ 9620] = 0;
        memory[ 9621] = 0;
        memory[ 9622] = 0;
        memory[ 9623] = 0;
        memory[ 9624] = 0;
        memory[ 9625] = 0;
        memory[ 9626] = 0;
        memory[ 9627] = 0;
        memory[ 9628] = 0;
        memory[ 9629] = 1;
        memory[ 9630] = 0;
        memory[ 9631] = 0;
        memory[ 9632] = 0;
        memory[ 9633] = 0;
        memory[ 9634] = 0;
        memory[ 9635] = 0;
        memory[ 9636] = 0;
        memory[ 9637] = 1;
        memory[ 9638] = 0;
        memory[ 9639] = 1;
        memory[ 9640] = 0;
        memory[ 9641] = 0;
        memory[ 9642] = 0;
        memory[ 9643] = 0;
        memory[ 9644] = 0;
        memory[ 9645] = 1;
        memory[ 9646] = 0;
        memory[ 9647] = 0;
        memory[ 9648] = 0;
        memory[ 9649] = 0;
        memory[ 9650] = 0;
        memory[ 9651] = 0;
        memory[ 9652] = 0;
        memory[ 9653] = 0;
        memory[ 9654] = 0;
        memory[ 9655] = 0;
        memory[ 9656] = 0;
        memory[ 9657] = 0;
        memory[ 9658] = 0;
        memory[ 9659] = 0;
        memory[ 9660] = 0;
        memory[ 9661] = 0;
        memory[ 9662] = 0;
        memory[ 9663] = 0;
        memory[ 9664] = 0;
        memory[ 9665] = 0;
        memory[ 9666] = 0;
        memory[ 9667] = 0;
        memory[ 9668] = 0;
        memory[ 9669] = 0;
        memory[ 9670] = 0;
        memory[ 9671] = 0;
        memory[ 9672] = 1;
        memory[ 9673] = 0;
        memory[ 9674] = 0;
        memory[ 9675] = 0;
        memory[ 9676] = 1;
        memory[ 9677] = 0;
        memory[ 9678] = 0;
        memory[ 9679] = 0;
        memory[ 9680] = 0;
        memory[ 9681] = 0;
        memory[ 9682] = 0;
        memory[ 9683] = 0;
        memory[ 9684] = 0;
        memory[ 9685] = 0;
        memory[ 9686] = 0;
        memory[ 9687] = 0;
        memory[ 9688] = 0;
        memory[ 9689] = 0;
        memory[ 9690] = 0;
        memory[ 9691] = 0;
        memory[ 9692] = 0;
        memory[ 9693] = 0;
        memory[ 9694] = 0;
        memory[ 9695] = 0;
        memory[ 9696] = 0;
        memory[ 9697] = 1;
        memory[ 9698] = 1;
        memory[ 9699] = 0;
        memory[ 9700] = 1;
        memory[ 9701] = 0;
        memory[ 9702] = 0;
        memory[ 9703] = 0;
        memory[ 9704] = 1;
        memory[ 9705] = 1;
        memory[ 9706] = 1;
        memory[ 9707] = 0;
        memory[ 9708] = 0;
        memory[ 9709] = 0;
        memory[ 9710] = 0;
        memory[ 9711] = 1;
        memory[ 9712] = 0;
        memory[ 9713] = 0;
        memory[ 9714] = 0;
        memory[ 9715] = 0;
        memory[ 9716] = 0;
        memory[ 9717] = 0;
        memory[ 9718] = 0;
        memory[ 9719] = 0;
        memory[ 9720] = 0;
        memory[ 9721] = 0;
        memory[ 9722] = 0;
        memory[ 9723] = 0;
        memory[ 9724] = 1;
        memory[ 9725] = 1;
        memory[ 9726] = 0;
        memory[ 9727] = 0;
        memory[ 9728] = 0;
        memory[ 9729] = 0;
        memory[ 9730] = 0;
        memory[ 9731] = 0;
        memory[ 9732] = 1;
        memory[ 9733] = 1;
        memory[ 9734] = 0;
        memory[ 9735] = 0;
        memory[ 9736] = 0;
        memory[ 9737] = 0;
        memory[ 9738] = 0;
        memory[ 9739] = 0;
        memory[ 9740] = 0;
        memory[ 9741] = 0;
        memory[ 9742] = 0;
        memory[ 9743] = 0;
        memory[ 9744] = 0;
        memory[ 9745] = 0;
        memory[ 9746] = 0;
        memory[ 9747] = 0;
        memory[ 9748] = 0;
        memory[ 9749] = 0;
        memory[ 9750] = 0;
        memory[ 9751] = 0;
        memory[ 9752] = 0;
        memory[ 9753] = 0;
        memory[ 9754] = 0;
        memory[ 9755] = 0;
        memory[ 9756] = 0;
        memory[ 9757] = 0;
        memory[ 9758] = 0;
        memory[ 9759] = 0;
        memory[ 9760] = 1;
        memory[ 9761] = 0;
        memory[ 9762] = 0;
        memory[ 9763] = 0;
        memory[ 9764] = 1;
        memory[ 9765] = 0;
        memory[ 9766] = 0;
        memory[ 9767] = 0;
        memory[ 9768] = 0;
        memory[ 9769] = 0;
        memory[ 9770] = 0;
        memory[ 9771] = 0;
        memory[ 9772] = 0;
        memory[ 9773] = 0;
        memory[ 9774] = 0;
        memory[ 9775] = 0;
        memory[ 9776] = 0;
        memory[ 9777] = 0;
        memory[ 9778] = 0;
        memory[ 9779] = 0;
        memory[ 9780] = 1;
        memory[ 9781] = 1;
        memory[ 9782] = 0;
        memory[ 9783] = 0;
        memory[ 9784] = 0;
        memory[ 9785] = 0;
        memory[ 9786] = 0;
        memory[ 9787] = 0;
        memory[ 9788] = 1;
        memory[ 9789] = 1;
        memory[ 9790] = 0;
        memory[ 9791] = 0;
        memory[ 9792] = 0;
        memory[ 9793] = 0;
        memory[ 9794] = 0;
        memory[ 9795] = 0;
        memory[ 9796] = 0;
        memory[ 9797] = 0;
        memory[ 9798] = 0;
        memory[ 9799] = 1;
        memory[ 9800] = 0;
        memory[ 9801] = 0;
        memory[ 9802] = 0;
        memory[ 9803] = 0;
        memory[ 9804] = 0;
        memory[ 9805] = 0;
        memory[ 9806] = 1;
        memory[ 9807] = 1;
        memory[ 9808] = 1;
        memory[ 9809] = 0;
        memory[ 9810] = 0;
        memory[ 9811] = 0;
        memory[ 9812] = 0;
        memory[ 9813] = 0;
        memory[ 9814] = 0;
        memory[ 9815] = 1;
        memory[ 9816] = 0;
        memory[ 9817] = 0;
        memory[ 9818] = 0;
        memory[ 9819] = 0;
        memory[ 9820] = 1;
        memory[ 9821] = 1;
        memory[ 9822] = 0;
        memory[ 9823] = 0;
        memory[ 9824] = 0;
        memory[ 9825] = 0;
        memory[ 9826] = 0;
        memory[ 9827] = 1;
        memory[ 9828] = 1;
        memory[ 9829] = 0;
        memory[ 9830] = 0;
        memory[ 9831] = 0;
        memory[ 9832] = 0;
        memory[ 9833] = 0;
        memory[ 9834] = 0;
        memory[ 9835] = 0;
        memory[ 9836] = 0;
        memory[ 9837] = 0;
        memory[ 9838] = 0;
        memory[ 9839] = 1;
        memory[ 9840] = 0;
        memory[ 9841] = 0;
        memory[ 9842] = 1;
        memory[ 9843] = 0;
        memory[ 9844] = 0;
        memory[ 9845] = 0;
        memory[ 9846] = 0;
        memory[ 9847] = 0;
        memory[ 9848] = 0;
        memory[ 9849] = 0;
        memory[ 9850] = 0;
        memory[ 9851] = 0;
        memory[ 9852] = 0;
        memory[ 9853] = 0;
        memory[ 9854] = 0;
        memory[ 9855] = 0;
        memory[ 9856] = 0;
        memory[ 9857] = 0;
        memory[ 9858] = 0;
        memory[ 9859] = 0;
        memory[ 9860] = 0;
        memory[ 9861] = 0;
        memory[ 9862] = 0;
        memory[ 9863] = 1;
        memory[ 9864] = 1;
        memory[ 9865] = 0;
        memory[ 9866] = 0;
        memory[ 9867] = 0;
        memory[ 9868] = 0;
        memory[ 9869] = 0;
        memory[ 9870] = 0;
        memory[ 9871] = 0;
        memory[ 9872] = 0;
        memory[ 9873] = 0;
        memory[ 9874] = 0;
        memory[ 9875] = 0;
        memory[ 9876] = 0;
        memory[ 9877] = 0;
        memory[ 9878] = 0;
        memory[ 9879] = 0;
        memory[ 9880] = 0;
        memory[ 9881] = 0;
        memory[ 9882] = 0;
        memory[ 9883] = 0;
        memory[ 9884] = 1;
        memory[ 9885] = 0;
        memory[ 9886] = 0;
        memory[ 9887] = 0;
        memory[ 9888] = 0;
        memory[ 9889] = 0;
        memory[ 9890] = 0;
        memory[ 9891] = 0;
        memory[ 9892] = 0;
        memory[ 9893] = 0;
        memory[ 9894] = 1;
        memory[ 9895] = 1;
        memory[ 9896] = 0;
        memory[ 9897] = 0;
        memory[ 9898] = 0;
        memory[ 9899] = 0;
        memory[ 9900] = 0;
        memory[ 9901] = 0;
        memory[ 9902] = 0;
        memory[ 9903] = 0;
        memory[ 9904] = 0;
        memory[ 9905] = 0;
        memory[ 9906] = 0;
        memory[ 9907] = 0;
        memory[ 9908] = 1;
        memory[ 9909] = 0;
        memory[ 9910] = 0;
        memory[ 9911] = 0;
        memory[ 9912] = 0;
        memory[ 9913] = 0;
        memory[ 9914] = 0;
        memory[ 9915] = 0;
        memory[ 9916] = 0;
        memory[ 9917] = 0;
        memory[ 9918] = 0;
        memory[ 9919] = 0;
        memory[ 9920] = 0;
        memory[ 9921] = 0;
        memory[ 9922] = 0;
        memory[ 9923] = 0;
        memory[ 9924] = 0;
        memory[ 9925] = 0;
        memory[ 9926] = 0;
        memory[ 9927] = 0;
        memory[ 9928] = 0;
        memory[ 9929] = 0;
        memory[ 9930] = 0;
        memory[ 9931] = 0;
        memory[ 9932] = 0;
        memory[ 9933] = 0;
        memory[ 9934] = 0;
        memory[ 9935] = 0;
        memory[ 9936] = 0;
        memory[ 9937] = 0;
        memory[ 9938] = 1;
        memory[ 9939] = 0;
        memory[ 9940] = 0;
        memory[ 9941] = 0;
        memory[ 9942] = 0;
        memory[ 9943] = 0;
        memory[ 9944] = 0;
        memory[ 9945] = 0;
        memory[ 9946] = 0;
        memory[ 9947] = 0;
        memory[ 9948] = 0;
        memory[ 9949] = 0;
        memory[ 9950] = 0;
        memory[ 9951] = 0;
        memory[ 9952] = 0;
        memory[ 9953] = 0;
        memory[ 9954] = 1;
        memory[ 9955] = 0;
        memory[ 9956] = 0;
        memory[ 9957] = 0;
        memory[ 9958] = 0;
        memory[ 9959] = 0;
        memory[ 9960] = 1;
        memory[ 9961] = 1;
        memory[ 9962] = 0;
        memory[ 9963] = 0;
        memory[ 9964] = 0;
        memory[ 9965] = 0;
        memory[ 9966] = 0;
        memory[ 9967] = 0;
        memory[ 9968] = 0;
        memory[ 9969] = 0;
        memory[ 9970] = 0;
        memory[ 9971] = 0;
        memory[ 9972] = 0;
        memory[ 9973] = 0;
        memory[ 9974] = 0;
        memory[ 9975] = 1;
        memory[ 9976] = 1;
        memory[ 9977] = 1;
        memory[ 9978] = 0;
        memory[ 9979] = 0;
        memory[ 9980] = 0;
        memory[ 9981] = 0;
        memory[ 9982] = 0;
        memory[ 9983] = 0;
        memory[ 9984] = 0;
        memory[ 9985] = 0;
        memory[ 9986] = 1;
        memory[ 9987] = 1;
        memory[ 9988] = 0;
        memory[ 9989] = 0;
        memory[ 9990] = 0;
        memory[ 9991] = 1;
        memory[ 9992] = 0;
        memory[ 9993] = 0;
        memory[ 9994] = 0;
        memory[ 9995] = 0;
        memory[ 9996] = 0;
        memory[ 9997] = 0;
        memory[ 9998] = 0;
        memory[ 9999] = 0;
        memory[10000] = 1;
        memory[10001] = 0;
        memory[10002] = 0;
        memory[10003] = 0;
        memory[10004] = 0;
        memory[10005] = 0;
        memory[10006] = 0;
        memory[10007] = 0;
        memory[10008] = 0;
        memory[10009] = 0;
        memory[10010] = 0;
        memory[10011] = 0;
        memory[10012] = 0;
        memory[10013] = 0;
        memory[10014] = 0;
        memory[10015] = 0;
        memory[10016] = 0;
        memory[10017] = 0;
        memory[10018] = 1;
        memory[10019] = 1;
        memory[10020] = 0;
        memory[10021] = 1;
        memory[10022] = 1;
        memory[10023] = 0;
        memory[10024] = 0;
        memory[10025] = 0;
        memory[10026] = 0;
        memory[10027] = 0;
        memory[10028] = 0;
        memory[10029] = 0;
        memory[10030] = 0;
        memory[10031] = 0;
        memory[10032] = 0;
        memory[10033] = 0;
        memory[10034] = 0;
        memory[10035] = 0;
        memory[10036] = 0;
        memory[10037] = 0;
        memory[10038] = 0;
        memory[10039] = 0;
        memory[10040] = 0;
        memory[10041] = 0;
        memory[10042] = 0;
        memory[10043] = 0;
        memory[10044] = 0;
        memory[10045] = 1;
        memory[10046] = 1;
        memory[10047] = 0;
        memory[10048] = 0;
        memory[10049] = 0;
        memory[10050] = 0;
        memory[10051] = 0;
        memory[10052] = 0;
        memory[10053] = 1;
        memory[10054] = 1;
        memory[10055] = 0;
        memory[10056] = 0;
        memory[10057] = 0;
        memory[10058] = 0;
        memory[10059] = 0;
        memory[10060] = 0;
        memory[10061] = 0;
        memory[10062] = 0;
        memory[10063] = 0;
        memory[10064] = 0;
        memory[10065] = 0;
        memory[10066] = 0;
        memory[10067] = 0;
        memory[10068] = 0;
        memory[10069] = 0;
        memory[10070] = 0;
        memory[10071] = 0;
        memory[10072] = 0;
        memory[10073] = 0;
        memory[10074] = 0;
        memory[10075] = 0;
        memory[10076] = 0;
        memory[10077] = 1;
        memory[10078] = 0;
        memory[10079] = 0;
        memory[10080] = 0;
        memory[10081] = 0;
        memory[10082] = 0;
        memory[10083] = 0;
        memory[10084] = 0;
        memory[10085] = 1;
        memory[10086] = 0;
        memory[10087] = 0;
        memory[10088] = 0;
        memory[10089] = 1;
        memory[10090] = 0;
        memory[10091] = 0;
        memory[10092] = 0;
        memory[10093] = 0;
        memory[10094] = 0;
        memory[10095] = 0;
        memory[10096] = 0;
        memory[10097] = 0;
        memory[10098] = 0;
        memory[10099] = 0;
        memory[10100] = 0;
        memory[10101] = 0;
        memory[10102] = 0;
        memory[10103] = 0;
        memory[10104] = 0;
        memory[10105] = 0;
        memory[10106] = 0;
        memory[10107] = 0;
        memory[10108] = 1;
        memory[10109] = 0;
        memory[10110] = 0;
        memory[10111] = 1;
        memory[10112] = 0;
        memory[10113] = 0;
        memory[10114] = 0;
        memory[10115] = 0;
        memory[10116] = 0;
        memory[10117] = 0;
        memory[10118] = 0;
        memory[10119] = 0;
        memory[10120] = 0;
        memory[10121] = 0;
        memory[10122] = 0;
        memory[10123] = 0;
        memory[10124] = 0;
        memory[10125] = 1;
        memory[10126] = 0;
        memory[10127] = 0;
        memory[10128] = 0;
        memory[10129] = 0;
        memory[10130] = 0;
        memory[10131] = 0;
        memory[10132] = 0;
        memory[10133] = 0;
        memory[10134] = 0;
        memory[10135] = 0;
        memory[10136] = 0;
        memory[10137] = 0;
        memory[10138] = 0;
        memory[10139] = 0;
        memory[10140] = 0;
        memory[10141] = 0;
        memory[10142] = 0;
        memory[10143] = 0;
        memory[10144] = 0;
        memory[10145] = 0;
        memory[10146] = 0;
        memory[10147] = 0;
        memory[10148] = 0;
        memory[10149] = 1;
        memory[10150] = 1;
        memory[10151] = 1;
        memory[10152] = 1;
        memory[10153] = 0;
        memory[10154] = 0;
        memory[10155] = 0;
        memory[10156] = 0;
        memory[10157] = 0;
        memory[10158] = 0;
        memory[10159] = 0;
        memory[10160] = 0;
        memory[10161] = 0;
        memory[10162] = 0;
        memory[10163] = 0;
        memory[10164] = 0;
        memory[10165] = 0;
        memory[10166] = 0;
        memory[10167] = 0;
        memory[10168] = 1;
        memory[10169] = 0;
        memory[10170] = 0;
        memory[10171] = 0;
        memory[10172] = 0;
        memory[10173] = 0;
        memory[10174] = 0;
        memory[10175] = 0;
        memory[10176] = 0;
        memory[10177] = 0;
        memory[10178] = 1;
        memory[10179] = 0;
        memory[10180] = 0;
        memory[10181] = 1;
        memory[10182] = 1;
        memory[10183] = 0;
        memory[10184] = 0;
        memory[10185] = 0;
        memory[10186] = 1;
        memory[10187] = 0;
        memory[10188] = 0;
        memory[10189] = 0;
        memory[10190] = 1;
        memory[10191] = 0;
        memory[10192] = 0;
        memory[10193] = 0;
        memory[10194] = 0;
        memory[10195] = 0;
        memory[10196] = 0;
        memory[10197] = 0;
        memory[10198] = 1;
        memory[10199] = 0;
        memory[10200] = 0;
        memory[10201] = 0;
        memory[10202] = 0;
        memory[10203] = 0;
        memory[10204] = 0;
        memory[10205] = 0;
        memory[10206] = 0;
        memory[10207] = 0;
        memory[10208] = 0;
        memory[10209] = 0;
        memory[10210] = 0;
        memory[10211] = 0;
        memory[10212] = 0;
        memory[10213] = 0;
        memory[10214] = 0;
        memory[10215] = 0;
        memory[10216] = 1;
        memory[10217] = 0;
        memory[10218] = 0;
        memory[10219] = 0;
        memory[10220] = 0;
        memory[10221] = 0;
        memory[10222] = 0;
        memory[10223] = 0;
        memory[10224] = 0;
        memory[10225] = 0;
        memory[10226] = 0;
        memory[10227] = 0;
        memory[10228] = 1;
        memory[10229] = 0;
        memory[10230] = 0;
        memory[10231] = 0;
        memory[10232] = 0;
        memory[10233] = 0;
        memory[10234] = 0;
        memory[10235] = 0;
        memory[10236] = 0;
        memory[10237] = 0;
        memory[10238] = 1;
        memory[10239] = 0;
        memory[10240] = 0;
        memory[10241] = 0;
        memory[10242] = 0;
        memory[10243] = 0;
        memory[10244] = 0;
        memory[10245] = 0;
        memory[10246] = 0;
        memory[10247] = 0;
        memory[10248] = 0;
        memory[10249] = 1;
        memory[10250] = 0;
        memory[10251] = 0;
        memory[10252] = 0;
        memory[10253] = 0;
        memory[10254] = 0;
        memory[10255] = 0;
        memory[10256] = 0;
        memory[10257] = 0;
        memory[10258] = 0;
        memory[10259] = 0;
        memory[10260] = 0;
        memory[10261] = 0;
        memory[10262] = 0;
        memory[10263] = 0;
        memory[10264] = 0;
        memory[10265] = 1;
        memory[10266] = 0;
        memory[10267] = 0;
        memory[10268] = 0;
        memory[10269] = 0;
        memory[10270] = 0;
        memory[10271] = 0;
        memory[10272] = 0;
        memory[10273] = 1;
        memory[10274] = 0;
        memory[10275] = 0;
        memory[10276] = 0;
        memory[10277] = 0;
        memory[10278] = 0;
        memory[10279] = 0;
        memory[10280] = 0;
        memory[10281] = 0;
        memory[10282] = 0;
        memory[10283] = 0;
        memory[10284] = 0;
        memory[10285] = 0;
        memory[10286] = 0;
        memory[10287] = 0;
        memory[10288] = 0;
        memory[10289] = 0;
        memory[10290] = 0;
        memory[10291] = 0;
        memory[10292] = 1;
        memory[10293] = 0;
        memory[10294] = 0;
        memory[10295] = 0;
        memory[10296] = 0;
        memory[10297] = 0;
        memory[10298] = 0;
        memory[10299] = 0;
        memory[10300] = 0;
        memory[10301] = 0;
        memory[10302] = 0;
        memory[10303] = 0;
        memory[10304] = 0;
        memory[10305] = 0;
        memory[10306] = 0;
        memory[10307] = 0;
        memory[10308] = 0;
        memory[10309] = 0;
        memory[10310] = 0;
        memory[10311] = 0;
        memory[10312] = 0;
        memory[10313] = 0;
        memory[10314] = 1;
        memory[10315] = 0;
        memory[10316] = 0;
        memory[10317] = 0;
        memory[10318] = 0;
        memory[10319] = 0;
        memory[10320] = 1;
        memory[10321] = 0;
        memory[10322] = 0;
        memory[10323] = 0;
        memory[10324] = 0;
        memory[10325] = 0;
        memory[10326] = 0;
        memory[10327] = 0;
        memory[10328] = 0;
        memory[10329] = 0;
        memory[10330] = 1;
        memory[10331] = 0;
        memory[10332] = 0;
        memory[10333] = 0;
        memory[10334] = 0;
        memory[10335] = 0;
        memory[10336] = 0;
        memory[10337] = 0;
        memory[10338] = 0;
        memory[10339] = 0;
        memory[10340] = 0;
        memory[10341] = 1;
        memory[10342] = 0;
        memory[10343] = 0;
        memory[10344] = 0;
        memory[10345] = 0;
        memory[10346] = 0;
        memory[10347] = 0;
        memory[10348] = 0;
        memory[10349] = 0;
        memory[10350] = 0;
        memory[10351] = 1;
        memory[10352] = 0;
        memory[10353] = 0;
        memory[10354] = 0;
        memory[10355] = 0;
        memory[10356] = 0;
        memory[10357] = 0;
        memory[10358] = 0;
        memory[10359] = 0;
        memory[10360] = 0;
        memory[10361] = 0;
        memory[10362] = 1;
        memory[10363] = 1;
        memory[10364] = 1;
        memory[10365] = 1;
        memory[10366] = 0;
        memory[10367] = 0;
        memory[10368] = 0;
        memory[10369] = 1;
        memory[10370] = 1;
        memory[10371] = 0;
        memory[10372] = 0;
        memory[10373] = 0;
        memory[10374] = 0;
        memory[10375] = 0;
        memory[10376] = 0;
        memory[10377] = 0;
        memory[10378] = 0;
        memory[10379] = 0;
        memory[10380] = 0;
        memory[10381] = 0;
        memory[10382] = 0;
        memory[10383] = 0;
        memory[10384] = 0;
        memory[10385] = 0;
        memory[10386] = 0;
        memory[10387] = 0;
        memory[10388] = 0;
        memory[10389] = 0;
        memory[10390] = 0;
        memory[10391] = 0;
        memory[10392] = 0;
        memory[10393] = 0;
        memory[10394] = 0;
        memory[10395] = 0;
        memory[10396] = 0;
        memory[10397] = 0;
        memory[10398] = 0;
        memory[10399] = 0;
        memory[10400] = 0;
        memory[10401] = 0;
        memory[10402] = 0;
        memory[10403] = 0;
        memory[10404] = 0;
        memory[10405] = 0;
        memory[10406] = 0;
        memory[10407] = 0;
        memory[10408] = 1;
        memory[10409] = 1;
        memory[10410] = 0;
        memory[10411] = 0;
        memory[10412] = 0;
        memory[10413] = 0;
        memory[10414] = 0;
        memory[10415] = 0;
        memory[10416] = 0;
        memory[10417] = 0;
        memory[10418] = 0;
        memory[10419] = 0;
        memory[10420] = 0;
        memory[10421] = 0;
        memory[10422] = 0;
        memory[10423] = 0;
        memory[10424] = 0;
        memory[10425] = 0;
        memory[10426] = 0;
        memory[10427] = 0;
        memory[10428] = 1;
        memory[10429] = 0;
        memory[10430] = 0;
        memory[10431] = 0;
        memory[10432] = 0;
        memory[10433] = 0;
        memory[10434] = 0;
        memory[10435] = 0;
        memory[10436] = 1;
        memory[10437] = 0;
        memory[10438] = 0;
        memory[10439] = 0;
        memory[10440] = 1;
        memory[10441] = 0;
        memory[10442] = 0;
        memory[10443] = 0;
        memory[10444] = 0;
        memory[10445] = 0;
        memory[10446] = 0;
        memory[10447] = 0;
        memory[10448] = 0;
        memory[10449] = 0;
        memory[10450] = 0;
        memory[10451] = 0;
        memory[10452] = 0;
        memory[10453] = 0;
        memory[10454] = 0;
        memory[10455] = 0;
        memory[10456] = 0;
        memory[10457] = 0;
        memory[10458] = 0;
        memory[10459] = 0;
        memory[10460] = 0;
        memory[10461] = 0;
        memory[10462] = 0;
        memory[10463] = 0;
        memory[10464] = 0;
        memory[10465] = 0;
        memory[10466] = 1;
        memory[10467] = 1;
        memory[10468] = 0;
        memory[10469] = 0;
        memory[10470] = 0;
        memory[10471] = 0;
        memory[10472] = 0;
        memory[10473] = 0;
        memory[10474] = 0;
        memory[10475] = 0;
        memory[10476] = 0;
        memory[10477] = 0;
        memory[10478] = 0;
        memory[10479] = 0;
        memory[10480] = 0;
        memory[10481] = 0;
        memory[10482] = 0;
        memory[10483] = 0;
        memory[10484] = 0;
        memory[10485] = 0;
        memory[10486] = 0;
        memory[10487] = 0;
        memory[10488] = 0;
        memory[10489] = 0;
        memory[10490] = 0;
        memory[10491] = 0;
        memory[10492] = 1;
        memory[10493] = 0;
        memory[10494] = 0;
        memory[10495] = 0;
        memory[10496] = 0;
        memory[10497] = 0;
        memory[10498] = 0;
        memory[10499] = 0;
        memory[10500] = 0;
        memory[10501] = 0;
        memory[10502] = 0;
        memory[10503] = 0;
        memory[10504] = 0;
        memory[10505] = 0;
        memory[10506] = 0;
        memory[10507] = 0;
        memory[10508] = 0;
        memory[10509] = 0;
        memory[10510] = 1;
        memory[10511] = 0;
        memory[10512] = 0;
        memory[10513] = 0;
        memory[10514] = 0;
        memory[10515] = 0;
        memory[10516] = 0;
        memory[10517] = 0;
        memory[10518] = 0;
        memory[10519] = 0;
        memory[10520] = 0;
        memory[10521] = 0;
        memory[10522] = 0;
        memory[10523] = 0;
        memory[10524] = 0;
        memory[10525] = 0;
        memory[10526] = 0;
        memory[10527] = 1;
        memory[10528] = 0;
        memory[10529] = 0;
        memory[10530] = 0;
        memory[10531] = 0;
        memory[10532] = 0;
        memory[10533] = 0;
        memory[10534] = 0;
        memory[10535] = 0;
        memory[10536] = 0;
        memory[10537] = 0;
        memory[10538] = 0;
        memory[10539] = 0;
        memory[10540] = 1;
        memory[10541] = 0;
        memory[10542] = 0;
        memory[10543] = 0;
        memory[10544] = 1;
        memory[10545] = 0;
        memory[10546] = 0;
        memory[10547] = 0;
        memory[10548] = 0;
        memory[10549] = 0;
        memory[10550] = 0;
        memory[10551] = 1;
        memory[10552] = 1;
        memory[10553] = 1;
        memory[10554] = 1;
        memory[10555] = 0;
        memory[10556] = 0;
        memory[10557] = 0;
        memory[10558] = 0;
        memory[10559] = 0;
        memory[10560] = 0;
        memory[10561] = 0;
        memory[10562] = 0;
        memory[10563] = 1;
        memory[10564] = 0;
        memory[10565] = 0;
        memory[10566] = 0;
        memory[10567] = 0;
        memory[10568] = 0;
        memory[10569] = 0;
        memory[10570] = 0;
        memory[10571] = 0;
        memory[10572] = 0;
        memory[10573] = 0;
        memory[10574] = 0;
        memory[10575] = 0;
        memory[10576] = 0;
        memory[10577] = 0;
        memory[10578] = 0;
        memory[10579] = 0;
        memory[10580] = 0;
        memory[10581] = 0;
        memory[10582] = 0;
        memory[10583] = 0;
        memory[10584] = 1;
        memory[10585] = 0;
        memory[10586] = 0;
        memory[10587] = 0;
        memory[10588] = 1;
        memory[10589] = 1;
        memory[10590] = 0;
        memory[10591] = 0;
        memory[10592] = 0;
        memory[10593] = 0;
        memory[10594] = 0;
        memory[10595] = 0;
        memory[10596] = 0;
        memory[10597] = 0;
        memory[10598] = 0;
        memory[10599] = 0;
        memory[10600] = 0;
        memory[10601] = 0;
        memory[10602] = 0;
        memory[10603] = 0;
        memory[10604] = 1;
        memory[10605] = 0;
        memory[10606] = 0;
        memory[10607] = 0;
        memory[10608] = 0;
        memory[10609] = 0;
        memory[10610] = 0;
        memory[10611] = 0;
        memory[10612] = 0;
        memory[10613] = 0;
        memory[10614] = 0;
        memory[10615] = 0;
        memory[10616] = 0;
        memory[10617] = 0;
        memory[10618] = 1;
        memory[10619] = 0;
        memory[10620] = 1;
        memory[10621] = 1;
        memory[10622] = 1;
        memory[10623] = 0;
        memory[10624] = 0;
        memory[10625] = 0;
        memory[10626] = 0;
        memory[10627] = 0;
        memory[10628] = 0;
        memory[10629] = 0;
        memory[10630] = 0;
        memory[10631] = 0;
        memory[10632] = 0;
        memory[10633] = 0;
        memory[10634] = 0;
        memory[10635] = 0;
        memory[10636] = 0;
        memory[10637] = 0;
        memory[10638] = 0;
        memory[10639] = 0;
        memory[10640] = 0;
        memory[10641] = 0;
        memory[10642] = 0;
        memory[10643] = 0;
        memory[10644] = 0;
        memory[10645] = 0;
        memory[10646] = 0;
        memory[10647] = 0;
        memory[10648] = 0;
        memory[10649] = 0;
        memory[10650] = 0;
        memory[10651] = 0;
        memory[10652] = 0;
        memory[10653] = 0;
        memory[10654] = 0;
        memory[10655] = 0;
        memory[10656] = 0;
        memory[10657] = 0;
        memory[10658] = 0;
        memory[10659] = 0;
        memory[10660] = 0;
        memory[10661] = 0;
        memory[10662] = 0;
        memory[10663] = 0;
        memory[10664] = 0;
        memory[10665] = 0;
        memory[10666] = 0;
        memory[10667] = 0;
        memory[10668] = 0;
        memory[10669] = 0;
        memory[10670] = 0;
        memory[10671] = 0;
        memory[10672] = 0;
        memory[10673] = 0;
        memory[10674] = 0;
        memory[10675] = 0;
        memory[10676] = 0;
        memory[10677] = 0;
        memory[10678] = 0;
        memory[10679] = 0;
        memory[10680] = 0;
        memory[10681] = 0;
        memory[10682] = 0;
        memory[10683] = 1;
        memory[10684] = 0;
        memory[10685] = 0;
        memory[10686] = 0;
        memory[10687] = 0;
        memory[10688] = 1;
        memory[10689] = 0;
        memory[10690] = 0;
        memory[10691] = 0;
        memory[10692] = 0;
        memory[10693] = 0;
        memory[10694] = 0;
        memory[10695] = 0;
        memory[10696] = 0;
        memory[10697] = 0;
        memory[10698] = 0;
        memory[10699] = 0;
        memory[10700] = 0;
        memory[10701] = 0;
        memory[10702] = 0;
        memory[10703] = 0;
        memory[10704] = 0;
        memory[10705] = 0;
        memory[10706] = 0;
        memory[10707] = 0;
        memory[10708] = 0;
        memory[10709] = 0;
        memory[10710] = 0;
        memory[10711] = 0;
        memory[10712] = 0;
        memory[10713] = 0;
        memory[10714] = 1;
        memory[10715] = 0;
        memory[10716] = 0;
        memory[10717] = 0;
        memory[10718] = 0;
        memory[10719] = 0;
        memory[10720] = 0;
        memory[10721] = 0;
        memory[10722] = 0;
        memory[10723] = 0;
        memory[10724] = 0;
        memory[10725] = 1;
        memory[10726] = 0;
        memory[10727] = 0;
        memory[10728] = 0;
        memory[10729] = 0;
        memory[10730] = 0;
        memory[10731] = 0;
        memory[10732] = 0;
        memory[10733] = 0;
        memory[10734] = 0;
        memory[10735] = 0;
        memory[10736] = 0;
        memory[10737] = 0;
        memory[10738] = 0;
        memory[10739] = 0;
        memory[10740] = 0;
        memory[10741] = 0;
        memory[10742] = 0;
        memory[10743] = 0;
        memory[10744] = 0;
        memory[10745] = 0;
        memory[10746] = 0;
        memory[10747] = 0;
        memory[10748] = 0;
        memory[10749] = 0;
        memory[10750] = 0;
        memory[10751] = 0;
        memory[10752] = 1;
        memory[10753] = 0;
        memory[10754] = 0;
        memory[10755] = 0;
        memory[10756] = 0;
        memory[10757] = 0;
        memory[10758] = 0;
        memory[10759] = 0;
        memory[10760] = 0;
        memory[10761] = 0;
        memory[10762] = 0;
        memory[10763] = 0;
        memory[10764] = 0;
        memory[10765] = 0;
        memory[10766] = 0;
        memory[10767] = 0;
        memory[10768] = 0;
        memory[10769] = 0;
        memory[10770] = 0;
        memory[10771] = 0;
        memory[10772] = 0;
        memory[10773] = 0;
        memory[10774] = 0;
        memory[10775] = 0;
        memory[10776] = 0;
        memory[10777] = 0;
        memory[10778] = 0;
        memory[10779] = 0;
        memory[10780] = 1;
        memory[10781] = 0;
        memory[10782] = 0;
        memory[10783] = 1;
        memory[10784] = 0;
        memory[10785] = 0;
        memory[10786] = 0;
        memory[10787] = 0;
        memory[10788] = 0;
        memory[10789] = 1;
        memory[10790] = 0;
        memory[10791] = 0;
        memory[10792] = 1;
        memory[10793] = 1;
        memory[10794] = 0;
        memory[10795] = 0;
        memory[10796] = 0;
        memory[10797] = 0;
        memory[10798] = 0;
        memory[10799] = 0;
        memory[10800] = 0;
        memory[10801] = 0;
        memory[10802] = 0;
        memory[10803] = 0;
        memory[10804] = 0;
        memory[10805] = 0;
        memory[10806] = 0;
        memory[10807] = 1;
        memory[10808] = 0;
        memory[10809] = 0;
        memory[10810] = 1;
        memory[10811] = 1;
        memory[10812] = 0;
        memory[10813] = 0;
        memory[10814] = 0;
        memory[10815] = 1;
        memory[10816] = 0;
        memory[10817] = 0;
        memory[10818] = 0;
        memory[10819] = 0;
        memory[10820] = 0;
        memory[10821] = 0;
        memory[10822] = 1;
        memory[10823] = 0;
        memory[10824] = 0;
        memory[10825] = 0;
        memory[10826] = 0;
        memory[10827] = 0;
        memory[10828] = 0;
        memory[10829] = 0;
        memory[10830] = 0;
        memory[10831] = 0;
        memory[10832] = 0;
        memory[10833] = 1;
        memory[10834] = 1;
        memory[10835] = 0;
        memory[10836] = 0;
        memory[10837] = 0;
        memory[10838] = 0;
        memory[10839] = 0;
        memory[10840] = 0;
        memory[10841] = 0;
        memory[10842] = 0;
        memory[10843] = 0;
        memory[10844] = 0;
        memory[10845] = 0;
        memory[10846] = 1;
        memory[10847] = 0;
        memory[10848] = 0;
        memory[10849] = 0;
        memory[10850] = 0;
        memory[10851] = 0;
        memory[10852] = 0;
        memory[10853] = 0;
        memory[10854] = 0;
        memory[10855] = 0;
        memory[10856] = 0;
        memory[10857] = 0;
        memory[10858] = 0;
        memory[10859] = 0;
        memory[10860] = 0;
        memory[10861] = 0;
        memory[10862] = 0;
        memory[10863] = 0;
        memory[10864] = 0;
        memory[10865] = 0;
        memory[10866] = 0;
        memory[10867] = 0;
        memory[10868] = 0;
        memory[10869] = 0;
        memory[10870] = 0;
        memory[10871] = 0;
        memory[10872] = 0;
        memory[10873] = 0;
        memory[10874] = 0;
        memory[10875] = 0;
        memory[10876] = 0;
        memory[10877] = 0;
        memory[10878] = 0;
        memory[10879] = 0;
        memory[10880] = 0;
        memory[10881] = 0;
        memory[10882] = 0;
        memory[10883] = 0;
        memory[10884] = 0;
        memory[10885] = 0;
        memory[10886] = 0;
        memory[10887] = 1;
        memory[10888] = 0;
        memory[10889] = 1;
        memory[10890] = 0;
        memory[10891] = 0;
        memory[10892] = 0;
        memory[10893] = 0;
        memory[10894] = 0;
        memory[10895] = 0;
        memory[10896] = 0;
        memory[10897] = 0;
        memory[10898] = 0;
        memory[10899] = 1;
        memory[10900] = 0;
        memory[10901] = 0;
        memory[10902] = 0;
        memory[10903] = 0;
        memory[10904] = 0;
        memory[10905] = 0;
        memory[10906] = 1;
        memory[10907] = 0;
        memory[10908] = 0;
        memory[10909] = 0;
        memory[10910] = 0;
        memory[10911] = 0;
        memory[10912] = 1;
        memory[10913] = 0;
        memory[10914] = 0;
        memory[10915] = 0;
        memory[10916] = 0;
        memory[10917] = 1;
        memory[10918] = 0;
        memory[10919] = 0;
        memory[10920] = 0;
        memory[10921] = 0;
        memory[10922] = 1;
        memory[10923] = 0;
        memory[10924] = 0;
        memory[10925] = 0;
        memory[10926] = 0;
        memory[10927] = 0;
        memory[10928] = 0;
        memory[10929] = 0;
        memory[10930] = 0;
        memory[10931] = 0;
        memory[10932] = 0;
        memory[10933] = 0;
        memory[10934] = 0;
        memory[10935] = 0;
        memory[10936] = 0;
        memory[10937] = 0;
        memory[10938] = 0;
        memory[10939] = 0;
        memory[10940] = 0;
        memory[10941] = 0;
        memory[10942] = 0;
        memory[10943] = 0;
        memory[10944] = 0;
        memory[10945] = 0;
        memory[10946] = 0;
        memory[10947] = 0;
        memory[10948] = 0;
        memory[10949] = 0;
        memory[10950] = 0;
        memory[10951] = 0;
        memory[10952] = 0;
        memory[10953] = 0;
        memory[10954] = 0;
        memory[10955] = 0;
        memory[10956] = 1;
        memory[10957] = 0;
        memory[10958] = 0;
        memory[10959] = 1;
        memory[10960] = 0;
        memory[10961] = 0;
        memory[10962] = 0;
        memory[10963] = 0;
        memory[10964] = 0;
        memory[10965] = 0;
        memory[10966] = 1;
        memory[10967] = 0;
        memory[10968] = 0;
        memory[10969] = 0;
        memory[10970] = 0;
        memory[10971] = 0;
        memory[10972] = 0;
        memory[10973] = 0;
        memory[10974] = 0;
        memory[10975] = 0;
        memory[10976] = 0;
        memory[10977] = 0;
        memory[10978] = 1;
        memory[10979] = 0;
        memory[10980] = 0;
        memory[10981] = 0;
        memory[10982] = 0;
        memory[10983] = 0;
        memory[10984] = 0;
        memory[10985] = 0;
        memory[10986] = 0;
        memory[10987] = 0;
        memory[10988] = 1;
        memory[10989] = 1;
        memory[10990] = 0;
        memory[10991] = 0;
        memory[10992] = 0;
        memory[10993] = 0;
        memory[10994] = 0;
        memory[10995] = 0;
        memory[10996] = 1;
        memory[10997] = 1;
        memory[10998] = 0;
        memory[10999] = 0;
        memory[11000] = 0;
        memory[11001] = 0;
        memory[11002] = 0;
        memory[11003] = 0;
        memory[11004] = 1;
        memory[11005] = 0;
        memory[11006] = 0;
        memory[11007] = 0;
        memory[11008] = 0;
        memory[11009] = 0;
        memory[11010] = 0;
        memory[11011] = 0;
        memory[11012] = 0;
        memory[11013] = 0;
        memory[11014] = 0;
        memory[11015] = 0;
        memory[11016] = 1;
        memory[11017] = 0;
        memory[11018] = 0;
        memory[11019] = 0;
        memory[11020] = 0;
        memory[11021] = 1;
        memory[11022] = 1;
        memory[11023] = 0;
        memory[11024] = 0;
        memory[11025] = 0;
        memory[11026] = 0;
        memory[11027] = 0;
        memory[11028] = 0;
        memory[11029] = 0;
        memory[11030] = 0;
        memory[11031] = 1;
        memory[11032] = 0;
        memory[11033] = 0;
        memory[11034] = 0;
        memory[11035] = 0;
        memory[11036] = 0;
        memory[11037] = 0;
        memory[11038] = 0;
        memory[11039] = 0;
        memory[11040] = 0;
        memory[11041] = 0;
        memory[11042] = 0;
        memory[11043] = 0;
        memory[11044] = 0;
        memory[11045] = 0;
        memory[11046] = 1;
        memory[11047] = 0;
        memory[11048] = 0;
        memory[11049] = 0;
        memory[11050] = 0;
        memory[11051] = 0;
        memory[11052] = 0;
        memory[11053] = 0;
        memory[11054] = 0;
        memory[11055] = 0;
        memory[11056] = 0;
        memory[11057] = 0;
        memory[11058] = 0;
        memory[11059] = 0;
        memory[11060] = 0;
        memory[11061] = 0;
        memory[11062] = 0;
        memory[11063] = 1;
        memory[11064] = 0;
        memory[11065] = 0;
        memory[11066] = 0;
        memory[11067] = 0;
        memory[11068] = 0;
        memory[11069] = 0;
        memory[11070] = 0;
        memory[11071] = 0;
        memory[11072] = 0;
        memory[11073] = 0;
        memory[11074] = 0;
        memory[11075] = 0;
        memory[11076] = 1;
        memory[11077] = 0;
        memory[11078] = 0;
        memory[11079] = 0;
        memory[11080] = 0;
        memory[11081] = 1;
        memory[11082] = 0;
        memory[11083] = 0;
        memory[11084] = 0;
        memory[11085] = 0;
        memory[11086] = 0;
        memory[11087] = 0;
        memory[11088] = 0;
        memory[11089] = 0;
        memory[11090] = 0;
        memory[11091] = 0;
        memory[11092] = 0;
        memory[11093] = 0;
        memory[11094] = 0;
        memory[11095] = 0;
        memory[11096] = 0;
        memory[11097] = 0;
        memory[11098] = 0;
        memory[11099] = 1;
        memory[11100] = 1;
        memory[11101] = 0;
        memory[11102] = 0;
        memory[11103] = 0;
        memory[11104] = 0;
        memory[11105] = 0;
        memory[11106] = 0;
        memory[11107] = 0;
        memory[11108] = 0;
        memory[11109] = 0;
        memory[11110] = 0;
        memory[11111] = 1;
        memory[11112] = 0;
        memory[11113] = 0;
        memory[11114] = 0;
        memory[11115] = 0;
        memory[11116] = 0;
        memory[11117] = 0;
        memory[11118] = 0;
        memory[11119] = 0;
        memory[11120] = 0;
        memory[11121] = 0;
        memory[11122] = 0;
        memory[11123] = 0;
        memory[11124] = 0;
        memory[11125] = 0;
        memory[11126] = 0;
        memory[11127] = 0;
        memory[11128] = 0;
        memory[11129] = 0;
        memory[11130] = 1;
        memory[11131] = 0;
        memory[11132] = 0;
        memory[11133] = 0;
        memory[11134] = 0;
        memory[11135] = 0;
        memory[11136] = 0;
        memory[11137] = 0;
        memory[11138] = 0;
        memory[11139] = 0;
        memory[11140] = 0;
        memory[11141] = 0;
        memory[11142] = 0;
        memory[11143] = 0;
        memory[11144] = 0;
        memory[11145] = 0;
        memory[11146] = 0;
        memory[11147] = 0;
        memory[11148] = 0;
        memory[11149] = 0;
        memory[11150] = 0;
        memory[11151] = 0;
        memory[11152] = 0;
        memory[11153] = 1;
        memory[11154] = 0;
        memory[11155] = 0;
        memory[11156] = 0;
        memory[11157] = 0;
        memory[11158] = 0;
        memory[11159] = 0;
        memory[11160] = 0;
        memory[11161] = 0;
        memory[11162] = 0;
        memory[11163] = 0;
        memory[11164] = 0;
        memory[11165] = 1;
        memory[11166] = 0;
        memory[11167] = 0;
        memory[11168] = 0;
        memory[11169] = 0;
        memory[11170] = 0;
        memory[11171] = 1;
        memory[11172] = 1;
        memory[11173] = 0;
        memory[11174] = 0;
        memory[11175] = 0;
        memory[11176] = 0;
        memory[11177] = 0;
        memory[11178] = 1;
        memory[11179] = 0;
        memory[11180] = 0;
        memory[11181] = 0;
        memory[11182] = 0;
        memory[11183] = 0;
        memory[11184] = 0;
        memory[11185] = 0;
        memory[11186] = 0;
        memory[11187] = 0;
        memory[11188] = 0;
        memory[11189] = 0;
        memory[11190] = 0;
        memory[11191] = 0;
        memory[11192] = 1;
        memory[11193] = 0;
        memory[11194] = 0;
        memory[11195] = 0;
        memory[11196] = 0;
        memory[11197] = 0;
        memory[11198] = 1;
        memory[11199] = 1;
        memory[11200] = 0;
        memory[11201] = 0;
        memory[11202] = 0;
        memory[11203] = 0;
        memory[11204] = 1;
        memory[11205] = 0;
        memory[11206] = 0;
        memory[11207] = 0;
        memory[11208] = 0;
        memory[11209] = 0;
        memory[11210] = 0;
        memory[11211] = 0;
        memory[11212] = 0;
        memory[11213] = 0;
        memory[11214] = 0;
        memory[11215] = 0;
        memory[11216] = 0;
        memory[11217] = 0;
        memory[11218] = 0;
        memory[11219] = 0;
        memory[11220] = 0;
        memory[11221] = 0;
        memory[11222] = 0;
        memory[11223] = 0;
        memory[11224] = 0;
        memory[11225] = 1;
        memory[11226] = 0;
        memory[11227] = 0;
        memory[11228] = 0;
        memory[11229] = 0;
        memory[11230] = 0;
        memory[11231] = 0;
        memory[11232] = 0;
        memory[11233] = 0;
        memory[11234] = 0;
        memory[11235] = 0;
        memory[11236] = 0;
        memory[11237] = 0;
        memory[11238] = 1;
        memory[11239] = 0;
        memory[11240] = 0;
        memory[11241] = 0;
        memory[11242] = 0;
        memory[11243] = 0;
        memory[11244] = 0;
        memory[11245] = 0;
        memory[11246] = 0;
        memory[11247] = 1;
        memory[11248] = 0;
        memory[11249] = 0;
        memory[11250] = 0;
        memory[11251] = 0;
        memory[11252] = 0;
        memory[11253] = 0;
        memory[11254] = 0;
        memory[11255] = 0;
        memory[11256] = 0;
        memory[11257] = 0;
        memory[11258] = 0;
        memory[11259] = 0;
        memory[11260] = 0;
        memory[11261] = 0;
        memory[11262] = 1;
        memory[11263] = 1;
        memory[11264] = 0;
        memory[11265] = 0;
        memory[11266] = 0;
        memory[11267] = 1;
        memory[11268] = 1;
        memory[11269] = 0;
        memory[11270] = 0;
        memory[11271] = 0;
        memory[11272] = 0;
        memory[11273] = 0;
        memory[11274] = 0;
        memory[11275] = 0;
        memory[11276] = 0;
        memory[11277] = 0;
        memory[11278] = 0;
        memory[11279] = 0;
        memory[11280] = 0;
        memory[11281] = 0;
        memory[11282] = 0;
        memory[11283] = 0;
        memory[11284] = 0;
        memory[11285] = 0;
        memory[11286] = 0;
        memory[11287] = 0;
        memory[11288] = 0;
        memory[11289] = 0;
        memory[11290] = 0;
        memory[11291] = 0;
        memory[11292] = 0;
        memory[11293] = 1;
        memory[11294] = 0;
        memory[11295] = 0;
        memory[11296] = 0;
        memory[11297] = 0;
        memory[11298] = 0;
        memory[11299] = 0;
        memory[11300] = 0;
        memory[11301] = 0;
        memory[11302] = 0;
        memory[11303] = 0;
        memory[11304] = 0;
        memory[11305] = 0;
        memory[11306] = 0;
        memory[11307] = 0;
        memory[11308] = 0;
        memory[11309] = 0;
        memory[11310] = 0;
        memory[11311] = 0;
        memory[11312] = 0;
        memory[11313] = 0;
        memory[11314] = 0;
        memory[11315] = 0;
        memory[11316] = 0;
        memory[11317] = 0;
        memory[11318] = 0;
        memory[11319] = 0;
        memory[11320] = 0;
        memory[11321] = 1;
        memory[11322] = 0;
        memory[11323] = 0;
        memory[11324] = 0;
        memory[11325] = 0;
        memory[11326] = 0;
        memory[11327] = 0;
        memory[11328] = 0;
        memory[11329] = 0;
        memory[11330] = 0;
        memory[11331] = 0;
        memory[11332] = 0;
        memory[11333] = 0;
        memory[11334] = 0;
        memory[11335] = 0;
        memory[11336] = 0;
        memory[11337] = 1;
        memory[11338] = 0;
        memory[11339] = 0;
        memory[11340] = 0;
        memory[11341] = 0;
        memory[11342] = 0;
        memory[11343] = 0;
        memory[11344] = 0;
        memory[11345] = 0;
        memory[11346] = 0;
        memory[11347] = 0;
        memory[11348] = 0;
        memory[11349] = 0;
        memory[11350] = 0;
        memory[11351] = 0;
        memory[11352] = 0;
        memory[11353] = 0;
        memory[11354] = 0;
        memory[11355] = 0;
        memory[11356] = 0;
        memory[11357] = 1;
        memory[11358] = 1;
        memory[11359] = 0;
        memory[11360] = 0;
        memory[11361] = 0;
        memory[11362] = 0;
        memory[11363] = 0;
        memory[11364] = 0;
        memory[11365] = 0;
        memory[11366] = 1;
        memory[11367] = 0;
        memory[11368] = 0;
        memory[11369] = 0;
        memory[11370] = 0;
        memory[11371] = 0;
        memory[11372] = 0;
        memory[11373] = 0;
        memory[11374] = 1;
        memory[11375] = 0;
        memory[11376] = 0;
        memory[11377] = 0;
        memory[11378] = 0;
        memory[11379] = 0;
        memory[11380] = 0;
        memory[11381] = 1;
        memory[11382] = 0;
        memory[11383] = 0;
        memory[11384] = 0;
        memory[11385] = 0;
        memory[11386] = 0;
        memory[11387] = 0;
        memory[11388] = 0;
        memory[11389] = 0;
        memory[11390] = 0;
        memory[11391] = 0;
        memory[11392] = 0;
        memory[11393] = 1;
        memory[11394] = 0;
        memory[11395] = 0;
        memory[11396] = 0;
        memory[11397] = 0;
        memory[11398] = 0;
        memory[11399] = 0;
        memory[11400] = 0;
        memory[11401] = 0;
        memory[11402] = 0;
        memory[11403] = 0;
        memory[11404] = 0;
        memory[11405] = 1;
        memory[11406] = 0;
        memory[11407] = 0;
        memory[11408] = 0;
        memory[11409] = 0;
        memory[11410] = 0;
        memory[11411] = 0;
        memory[11412] = 0;
        memory[11413] = 1;
        memory[11414] = 1;
        memory[11415] = 0;
        memory[11416] = 0;
        memory[11417] = 0;
        memory[11418] = 0;
        memory[11419] = 0;
        memory[11420] = 0;
        memory[11421] = 0;
        memory[11422] = 0;
        memory[11423] = 0;
        memory[11424] = 0;
        memory[11425] = 0;
        memory[11426] = 0;
        memory[11427] = 1;
        memory[11428] = 0;
        memory[11429] = 0;
        memory[11430] = 0;
        memory[11431] = 0;
        memory[11432] = 0;
        memory[11433] = 0;
        memory[11434] = 0;
        memory[11435] = 0;
        memory[11436] = 0;
        memory[11437] = 0;
        memory[11438] = 0;
        memory[11439] = 0;
        memory[11440] = 0;
        memory[11441] = 0;
        memory[11442] = 0;
        memory[11443] = 0;
        memory[11444] = 0;
        memory[11445] = 0;
        memory[11446] = 0;
        memory[11447] = 0;
        memory[11448] = 0;
        memory[11449] = 0;
        memory[11450] = 1;
        memory[11451] = 1;
        memory[11452] = 0;
        memory[11453] = 1;
        memory[11454] = 0;
        memory[11455] = 0;
        memory[11456] = 0;
        memory[11457] = 0;
        memory[11458] = 0;
        memory[11459] = 0;
        memory[11460] = 1;
        memory[11461] = 1;
        memory[11462] = 0;
        memory[11463] = 0;
        memory[11464] = 0;
        memory[11465] = 0;
        memory[11466] = 0;
        memory[11467] = 0;
        memory[11468] = 0;
        memory[11469] = 0;
        memory[11470] = 0;
        memory[11471] = 0;
        memory[11472] = 0;
        memory[11473] = 0;
        memory[11474] = 0;
        memory[11475] = 0;
        memory[11476] = 1;
        memory[11477] = 0;
        memory[11478] = 1;
        memory[11479] = 1;
        memory[11480] = 1;
        memory[11481] = 0;
        memory[11482] = 0;
        memory[11483] = 0;
        memory[11484] = 0;
        memory[11485] = 0;
        memory[11486] = 0;
        memory[11487] = 0;
        memory[11488] = 0;
        memory[11489] = 1;
        memory[11490] = 1;
        memory[11491] = 1;
        memory[11492] = 0;
        memory[11493] = 0;
        memory[11494] = 0;
        memory[11495] = 0;
        memory[11496] = 0;
        memory[11497] = 1;
        memory[11498] = 0;
        memory[11499] = 0;
        memory[11500] = 0;
        memory[11501] = 0;
        memory[11502] = 0;
        memory[11503] = 0;
        memory[11504] = 0;
        memory[11505] = 0;
        memory[11506] = 0;
        memory[11507] = 0;
        memory[11508] = 0;
        memory[11509] = 0;
        memory[11510] = 0;
        memory[11511] = 1;
        memory[11512] = 0;
        memory[11513] = 1;
        memory[11514] = 0;
        memory[11515] = 0;
        memory[11516] = 0;
        memory[11517] = 0;
        memory[11518] = 0;
        memory[11519] = 0;
        memory[11520] = 0;
        memory[11521] = 0;
        memory[11522] = 0;
        memory[11523] = 0;
        memory[11524] = 0;
        memory[11525] = 0;
        memory[11526] = 0;
        memory[11527] = 0;
        memory[11528] = 1;
        memory[11529] = 1;
        memory[11530] = 0;
        memory[11531] = 0;
        memory[11532] = 0;
        memory[11533] = 0;
        memory[11534] = 1;
        memory[11535] = 1;
        memory[11536] = 0;
        memory[11537] = 0;
        memory[11538] = 0;
        memory[11539] = 0;
        memory[11540] = 0;
        memory[11541] = 0;
        memory[11542] = 0;
        memory[11543] = 0;
        memory[11544] = 0;
        memory[11545] = 0;
        memory[11546] = 0;
        memory[11547] = 0;
        memory[11548] = 0;
        memory[11549] = 0;
        memory[11550] = 0;
        memory[11551] = 0;
        memory[11552] = 0;
        memory[11553] = 0;
        memory[11554] = 0;
        memory[11555] = 0;
        memory[11556] = 0;
        memory[11557] = 0;
        memory[11558] = 0;
        memory[11559] = 0;
        memory[11560] = 0;
        memory[11561] = 0;
        memory[11562] = 0;
        memory[11563] = 0;
        memory[11564] = 0;
        memory[11565] = 0;
        memory[11566] = 0;
        memory[11567] = 0;
        memory[11568] = 0;
        memory[11569] = 0;
        memory[11570] = 0;
        memory[11571] = 0;
        memory[11572] = 0;
        memory[11573] = 0;
        memory[11574] = 0;
        memory[11575] = 0;
        memory[11576] = 1;
        memory[11577] = 1;
        memory[11578] = 0;
        memory[11579] = 0;
        memory[11580] = 0;
        memory[11581] = 0;
        memory[11582] = 0;
        memory[11583] = 0;
        memory[11584] = 0;
        memory[11585] = 0;
        memory[11586] = 0;
        memory[11587] = 0;
        memory[11588] = 0;
        memory[11589] = 0;
        memory[11590] = 0;
        memory[11591] = 0;
        memory[11592] = 0;
        memory[11593] = 1;
        memory[11594] = 1;
        memory[11595] = 0;
        memory[11596] = 0;
        memory[11597] = 0;
        memory[11598] = 0;
        memory[11599] = 0;
        memory[11600] = 0;
        memory[11601] = 0;
        memory[11602] = 0;
        memory[11603] = 0;
        memory[11604] = 0;
        memory[11605] = 0;
        memory[11606] = 0;
        memory[11607] = 1;
        memory[11608] = 0;
        memory[11609] = 0;
        memory[11610] = 0;
        memory[11611] = 0;
        memory[11612] = 0;
        memory[11613] = 0;
        memory[11614] = 0;
        memory[11615] = 0;
        memory[11616] = 0;
        memory[11617] = 1;
        memory[11618] = 0;
        memory[11619] = 0;
        memory[11620] = 0;
        memory[11621] = 0;
        memory[11622] = 0;
        memory[11623] = 0;
        memory[11624] = 0;
        memory[11625] = 0;
        memory[11626] = 0;
        memory[11627] = 0;
        memory[11628] = 0;
        memory[11629] = 0;
        memory[11630] = 0;
        memory[11631] = 0;
        memory[11632] = 0;
        memory[11633] = 0;
        memory[11634] = 0;
        memory[11635] = 0;
        memory[11636] = 0;
        memory[11637] = 0;
        memory[11638] = 0;
        memory[11639] = 0;
        memory[11640] = 0;
        memory[11641] = 0;
        memory[11642] = 0;
        memory[11643] = 0;
        memory[11644] = 0;
        memory[11645] = 0;
        memory[11646] = 1;
        memory[11647] = 0;
        memory[11648] = 0;
        memory[11649] = 0;
        memory[11650] = 1;
        memory[11651] = 0;
        memory[11652] = 0;
        memory[11653] = 0;
        memory[11654] = 0;
        memory[11655] = 0;
        memory[11656] = 1;
        memory[11657] = 1;
        memory[11658] = 1;
        memory[11659] = 0;
        memory[11660] = 1;
        memory[11661] = 0;
        memory[11662] = 0;
        memory[11663] = 0;
        memory[11664] = 0;
        memory[11665] = 0;
        memory[11666] = 0;
        memory[11667] = 0;
        memory[11668] = 0;
        memory[11669] = 0;
        memory[11670] = 0;
        memory[11671] = 0;
        memory[11672] = 1;
        memory[11673] = 1;
        memory[11674] = 1;
        memory[11675] = 0;
        memory[11676] = 0;
        memory[11677] = 0;
        memory[11678] = 0;
        memory[11679] = 0;
        memory[11680] = 0;
        memory[11681] = 0;
        memory[11682] = 0;
        memory[11683] = 0;
        memory[11684] = 0;
        memory[11685] = 0;
        memory[11686] = 0;
        memory[11687] = 0;
        memory[11688] = 0;
        memory[11689] = 0;
        memory[11690] = 0;
        memory[11691] = 0;
        memory[11692] = 0;
        memory[11693] = 0;
        memory[11694] = 1;
        memory[11695] = 1;
        memory[11696] = 1;
        memory[11697] = 0;
        memory[11698] = 0;
        memory[11699] = 0;
        memory[11700] = 0;
        memory[11701] = 1;
        memory[11702] = 0;
        memory[11703] = 0;
        memory[11704] = 0;
        memory[11705] = 1;
        memory[11706] = 0;
        memory[11707] = 0;
        memory[11708] = 0;
        memory[11709] = 0;
        memory[11710] = 0;
        memory[11711] = 0;
        memory[11712] = 1;
        memory[11713] = 1;
        memory[11714] = 0;
        memory[11715] = 0;
        memory[11716] = 0;
        memory[11717] = 0;
        memory[11718] = 0;
        memory[11719] = 0;
        memory[11720] = 0;
        memory[11721] = 0;
        memory[11722] = 0;
        memory[11723] = 0;
        memory[11724] = 0;
        memory[11725] = 0;
        memory[11726] = 0;
        memory[11727] = 0;
        memory[11728] = 0;
        memory[11729] = 0;
        memory[11730] = 0;
        memory[11731] = 0;
        memory[11732] = 0;
        memory[11733] = 0;
        memory[11734] = 0;
        memory[11735] = 0;
        memory[11736] = 0;
        memory[11737] = 0;
        memory[11738] = 0;
        memory[11739] = 0;
        memory[11740] = 0;
        memory[11741] = 0;
        memory[11742] = 1;
        memory[11743] = 0;
        memory[11744] = 0;
        memory[11745] = 0;
        memory[11746] = 0;
        memory[11747] = 0;
        memory[11748] = 1;
        memory[11749] = 0;
        memory[11750] = 0;
        memory[11751] = 0;
        memory[11752] = 0;
        memory[11753] = 0;
        memory[11754] = 0;
        memory[11755] = 0;
        memory[11756] = 0;
        memory[11757] = 0;
        memory[11758] = 0;
        memory[11759] = 0;
        memory[11760] = 0;
        memory[11761] = 0;
        memory[11762] = 0;
        memory[11763] = 0;
        memory[11764] = 0;
        memory[11765] = 0;
        memory[11766] = 0;
        memory[11767] = 0;
        memory[11768] = 0;
        memory[11769] = 0;
        memory[11770] = 0;
        memory[11771] = 0;
        memory[11772] = 0;
        memory[11773] = 0;
        memory[11774] = 0;
        memory[11775] = 1;
        memory[11776] = 0;
        memory[11777] = 0;
        memory[11778] = 0;
        memory[11779] = 0;
        memory[11780] = 0;
        memory[11781] = 0;
        memory[11782] = 1;
        memory[11783] = 0;
        memory[11784] = 0;
        memory[11785] = 0;
        memory[11786] = 0;
        memory[11787] = 0;
        memory[11788] = 0;
        memory[11789] = 0;
        memory[11790] = 0;
        memory[11791] = 0;
        memory[11792] = 0;
        memory[11793] = 0;
        memory[11794] = 0;
        memory[11795] = 1;
        memory[11796] = 0;
        memory[11797] = 0;
        memory[11798] = 0;
        memory[11799] = 0;
        memory[11800] = 0;
        memory[11801] = 1;
        memory[11802] = 0;
        memory[11803] = 0;
        memory[11804] = 0;
        memory[11805] = 0;
        memory[11806] = 0;
        memory[11807] = 0;
        memory[11808] = 0;
        memory[11809] = 1;
        memory[11810] = 1;
        memory[11811] = 0;
        memory[11812] = 0;
        memory[11813] = 0;
        memory[11814] = 0;
        memory[11815] = 0;
        memory[11816] = 0;
        memory[11817] = 0;
        memory[11818] = 0;
        memory[11819] = 0;
        memory[11820] = 0;
        memory[11821] = 0;
        memory[11822] = 0;
        memory[11823] = 0;
        memory[11824] = 0;
        memory[11825] = 0;
        memory[11826] = 0;
        memory[11827] = 0;
        memory[11828] = 1;
        memory[11829] = 0;
        memory[11830] = 1;
        memory[11831] = 0;
        memory[11832] = 0;
        memory[11833] = 0;
        memory[11834] = 0;
        memory[11835] = 0;
        memory[11836] = 0;
        memory[11837] = 1;
        memory[11838] = 1;
        memory[11839] = 0;
        memory[11840] = 0;
        memory[11841] = 0;
        memory[11842] = 1;
        memory[11843] = 0;
        memory[11844] = 0;
        memory[11845] = 0;
        memory[11846] = 0;
        memory[11847] = 0;
        memory[11848] = 0;
        memory[11849] = 0;
        memory[11850] = 0;
        memory[11851] = 0;
        memory[11852] = 1;
        memory[11853] = 0;
        memory[11854] = 0;
        memory[11855] = 0;
        memory[11856] = 0;
        memory[11857] = 0;
        memory[11858] = 0;
        memory[11859] = 0;
        memory[11860] = 0;
        memory[11861] = 0;
        memory[11862] = 0;
        memory[11863] = 0;
        memory[11864] = 0;
        memory[11865] = 0;
        memory[11866] = 0;
        memory[11867] = 1;
        memory[11868] = 1;
        memory[11869] = 0;
        memory[11870] = 0;
        memory[11871] = 0;
        memory[11872] = 0;
        memory[11873] = 0;
        memory[11874] = 1;
        memory[11875] = 1;
        memory[11876] = 0;
        memory[11877] = 0;
        memory[11878] = 0;
        memory[11879] = 0;
        memory[11880] = 0;
        memory[11881] = 0;
        memory[11882] = 0;
        memory[11883] = 1;
        memory[11884] = 0;
        memory[11885] = 0;
        memory[11886] = 0;
        memory[11887] = 0;
        memory[11888] = 0;
        memory[11889] = 1;
        memory[11890] = 0;
        memory[11891] = 0;
        memory[11892] = 0;
        memory[11893] = 0;
        memory[11894] = 0;
        memory[11895] = 0;
        memory[11896] = 1;
        memory[11897] = 1;
        memory[11898] = 0;
        memory[11899] = 0;
        memory[11900] = 0;
        memory[11901] = 1;
        memory[11902] = 0;
        memory[11903] = 0;
        memory[11904] = 0;
        memory[11905] = 0;
        memory[11906] = 0;
        memory[11907] = 0;
        memory[11908] = 0;
        memory[11909] = 0;
        memory[11910] = 0;
        memory[11911] = 0;
        memory[11912] = 1;
        memory[11913] = 0;
        memory[11914] = 0;
        memory[11915] = 0;
        memory[11916] = 0;
        memory[11917] = 0;
        memory[11918] = 0;
        memory[11919] = 0;
        memory[11920] = 0;
        memory[11921] = 0;
        memory[11922] = 0;
        memory[11923] = 1;
        memory[11924] = 0;
        memory[11925] = 0;
        memory[11926] = 0;
        memory[11927] = 0;
        memory[11928] = 0;
        memory[11929] = 0;
        memory[11930] = 0;
        memory[11931] = 0;
        memory[11932] = 0;
        memory[11933] = 0;
        memory[11934] = 0;
        memory[11935] = 0;
        memory[11936] = 0;
        memory[11937] = 0;
        memory[11938] = 0;
        memory[11939] = 0;
        memory[11940] = 0;
        memory[11941] = 0;
        memory[11942] = 0;
        memory[11943] = 1;
        memory[11944] = 0;
        memory[11945] = 0;
        memory[11946] = 0;
        memory[11947] = 0;
        memory[11948] = 0;
        memory[11949] = 0;
        memory[11950] = 0;
        memory[11951] = 0;
        memory[11952] = 0;
        memory[11953] = 0;
        memory[11954] = 1;
        memory[11955] = 0;
        memory[11956] = 0;
        memory[11957] = 0;
        memory[11958] = 0;
        memory[11959] = 0;
        memory[11960] = 1;
        memory[11961] = 0;
        memory[11962] = 0;
        memory[11963] = 0;
        memory[11964] = 0;
        memory[11965] = 0;
        memory[11966] = 0;
        memory[11967] = 0;
        memory[11968] = 1;
        memory[11969] = 1;
        memory[11970] = 0;
        memory[11971] = 0;
        memory[11972] = 0;
        memory[11973] = 0;
        memory[11974] = 0;
        memory[11975] = 1;
        memory[11976] = 1;
        memory[11977] = 0;
        memory[11978] = 1;
        memory[11979] = 1;
        memory[11980] = 1;
        memory[11981] = 1;
        memory[11982] = 1;
        memory[11983] = 1;
        memory[11984] = 1;
        memory[11985] = 1;
        memory[11986] = 1;
        memory[11987] = 0;
        memory[11988] = 0;
        memory[11989] = 0;
        memory[11990] = 0;
        memory[11991] = 0;
        memory[11992] = 0;
        memory[11993] = 0;
        memory[11994] = 0;
        memory[11995] = 0;
        memory[11996] = 0;
        memory[11997] = 0;
        memory[11998] = 0;
        memory[11999] = 0;
        memory[12000] = 0;
        memory[12001] = 0;
        memory[12002] = 0;
        memory[12003] = 0;
        memory[12004] = 0;
        memory[12005] = 0;
        memory[12006] = 0;
        memory[12007] = 0;
        memory[12008] = 0;
        memory[12009] = 0;
        memory[12010] = 1;
        memory[12011] = 0;
        memory[12012] = 0;
        memory[12013] = 1;
        memory[12014] = 1;
        memory[12015] = 0;
        memory[12016] = 0;
        memory[12017] = 0;
        memory[12018] = 0;
        memory[12019] = 0;
        memory[12020] = 0;
        memory[12021] = 0;
        memory[12022] = 0;
        memory[12023] = 0;
        memory[12024] = 0;
        memory[12025] = 0;
        memory[12026] = 0;
        memory[12027] = 0;
        memory[12028] = 0;
        memory[12029] = 0;
        memory[12030] = 0;
        memory[12031] = 1;
        memory[12032] = 0;
        memory[12033] = 0;
        memory[12034] = 0;
        memory[12035] = 0;
        memory[12036] = 0;
        memory[12037] = 0;
        memory[12038] = 0;
        memory[12039] = 1;
        memory[12040] = 0;
        memory[12041] = 0;
        memory[12042] = 0;
        memory[12043] = 0;
        memory[12044] = 0;
        memory[12045] = 0;
        memory[12046] = 0;
        memory[12047] = 0;
        memory[12048] = 0;
        memory[12049] = 0;
        memory[12050] = 1;
        memory[12051] = 1;
        memory[12052] = 0;
        memory[12053] = 0;
        memory[12054] = 0;
        memory[12055] = 1;
        memory[12056] = 1;
        memory[12057] = 0;
        memory[12058] = 0;
        memory[12059] = 0;
        memory[12060] = 0;
        memory[12061] = 0;
        memory[12062] = 0;
        memory[12063] = 0;
        memory[12064] = 0;
        memory[12065] = 1;
        memory[12066] = 0;
        memory[12067] = 0;
        memory[12068] = 0;
        memory[12069] = 1;
        memory[12070] = 0;
        memory[12071] = 0;
        memory[12072] = 0;
        memory[12073] = 0;
        memory[12074] = 0;
        memory[12075] = 0;
        memory[12076] = 0;
        memory[12077] = 0;
        memory[12078] = 0;
        memory[12079] = 0;
        memory[12080] = 0;
        memory[12081] = 0;
        memory[12082] = 0;
        memory[12083] = 0;
        memory[12084] = 0;
        memory[12085] = 0;
        memory[12086] = 0;
        memory[12087] = 0;
        memory[12088] = 0;
        memory[12089] = 0;
        memory[12090] = 0;
        memory[12091] = 0;
        memory[12092] = 0;
        memory[12093] = 0;
        memory[12094] = 0;
        memory[12095] = 0;
        memory[12096] = 0;
        memory[12097] = 0;
        memory[12098] = 0;
        memory[12099] = 1;
        memory[12100] = 0;
        memory[12101] = 0;
        memory[12102] = 0;
        memory[12103] = 1;
        memory[12104] = 0;
        memory[12105] = 0;
        memory[12106] = 0;
        memory[12107] = 0;
        memory[12108] = 0;
        memory[12109] = 0;
        memory[12110] = 0;
        memory[12111] = 0;
        memory[12112] = 0;
        memory[12113] = 0;
        memory[12114] = 0;
        memory[12115] = 0;
        memory[12116] = 1;
        memory[12117] = 1;
        memory[12118] = 0;
        memory[12119] = 0;
        memory[12120] = 0;
        memory[12121] = 0;
        memory[12122] = 0;
        memory[12123] = 0;
        memory[12124] = 1;
        memory[12125] = 0;
        memory[12126] = 0;
        memory[12127] = 0;
        memory[12128] = 0;
        memory[12129] = 0;
        memory[12130] = 0;
        memory[12131] = 0;
        memory[12132] = 0;
        memory[12133] = 0;
        memory[12134] = 1;
        memory[12135] = 0;
        memory[12136] = 0;
        memory[12137] = 0;
        memory[12138] = 1;
        memory[12139] = 0;
        memory[12140] = 0;
        memory[12141] = 0;
        memory[12142] = 1;
        memory[12143] = 1;
        memory[12144] = 1;
        memory[12145] = 1;
        memory[12146] = 1;
        memory[12147] = 1;
        memory[12148] = 1;
        memory[12149] = 1;
        memory[12150] = 1;
        memory[12151] = 1;
        memory[12152] = 0;
        memory[12153] = 1;
        memory[12154] = 1;
        memory[12155] = 1;
        memory[12156] = 1;
        memory[12157] = 1;
        memory[12158] = 1;
        memory[12159] = 0;
        memory[12160] = 0;
        memory[12161] = 0;
        memory[12162] = 0;
        memory[12163] = 1;
        memory[12164] = 1;
        memory[12165] = 1;
        memory[12166] = 0;
        memory[12167] = 0;
        memory[12168] = 1;
        memory[12169] = 0;
        memory[12170] = 0;
        memory[12171] = 0;
        memory[12172] = 0;
        memory[12173] = 0;
        memory[12174] = 1;
        memory[12175] = 1;
        memory[12176] = 0;
        memory[12177] = 0;
        memory[12178] = 0;
        memory[12179] = 0;
        memory[12180] = 0;
        memory[12181] = 1;
        memory[12182] = 1;
        memory[12183] = 1;
        memory[12184] = 1;
        memory[12185] = 1;
        memory[12186] = 1;
        memory[12187] = 0;
        memory[12188] = 1;
        memory[12189] = 1;
        memory[12190] = 1;
        memory[12191] = 1;
        memory[12192] = 0;
        memory[12193] = 0;
        memory[12194] = 1;
        memory[12195] = 0;
        memory[12196] = 0;
        memory[12197] = 0;
        memory[12198] = 1;
        memory[12199] = 0;
        memory[12200] = 1;
        memory[12201] = 1;
        memory[12202] = 1;
        memory[12203] = 1;
        memory[12204] = 0;
        memory[12205] = 0;
        memory[12206] = 1;
        memory[12207] = 1;
        memory[12208] = 1;
        memory[12209] = 1;
        memory[12210] = 0;
        memory[12211] = 1;
        memory[12212] = 1;
        memory[12213] = 0;
        memory[12214] = 0;
        memory[12215] = 0;
        memory[12216] = 1;
        memory[12217] = 1;
        memory[12218] = 1;
        memory[12219] = 0;
        memory[12220] = 0;
        memory[12221] = 0;
        memory[12222] = 1;
        memory[12223] = 1;
    end

    always @(posedge clk) begin
        data <= memory[addr];
    end

endmodule
