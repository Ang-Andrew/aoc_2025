localparam NUM_NODES = 8;
localparam OUT_NODE = 0;
localparam YOU_NODE = 7;
