localparam WIDTH = 21;
localparam HEIGHT = 4;
localparam MEM_SIZE = 84;
