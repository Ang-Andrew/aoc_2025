localparam NUM_POINTS = 496;
