localparam WIDTH = 3725;
localparam HEIGHT = 5;
localparam COL_BITS = 40;
