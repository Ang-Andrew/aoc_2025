localparam WIDTH = 141;
localparam HEIGHT = 142;
localparam ROW_BITS = 282;
