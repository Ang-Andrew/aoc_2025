localparam NUM_NODES = 20;
localparam NUM_EDGES = 10;
localparam K_LIMIT = 10;
